----------------------------------------------------------------------------------
-- Company: Hatlab@Pitt
-- Author : Chao Zhou
-- Reference : 
-- Create Date: 07/25/2018
-- Description : Change the incoming signal into the form that is suitable for the Divison block(1.15 bit_shift, i.e. 1 integer 15 fractional bits). 
--               1)Use XOR gate to find the sign of result then convert the input to abs value
--               2)Find MSB and shift it to the first bit
--               3)Record the difference of number of bits shiffted for final reduction.
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use std.textio.all;


entity Div_Comb_Norm_tb is	
end Div_Comb_Norm_tb;

architecture Behavioral of Div_Comb_Norm_tb is

  constant c_clk_period  : time:=10 ns;
 
  
  signal r_N_in       : std_logic_vector(15 downto 0);
  signal r_D_in       : std_logic_vector(15 downto 0);
  signal w_sign       : std_logic :='0';
  signal w_bit_shift  : std_logic_vector(3 downto 0);
  signal w_N_out      : std_logic_vector(15 downto 0);
  signal w_D_out      : std_logic_vector(15 downto 0);
  signal w_Q_out      : std_logic_vector(15 downto 0);
  
  signal r_rst     : std_logic:='0';
  signal r_clk     : std_logic:='0';
  
  component Div_FormConv_Norm is
    port(
	N_in  : in std_logic_vector(15 downto 0);
	D_in  : in std_logic_vector(15 downto 0);   --Assume 16 bits income
	
	sign      : out std_logic := '0';
	bit_shift : out std_logic_vector (3 downto 0) := "0000";  --Also assume Denorminator is always graeator than Norminator
	
	N_out     : out std_logic_vector(15 downto 0):= (others => '1');
	D_out     : out std_logic_vector(15 downto 0):= (others => '1');
	
	clk : in std_logic;
	rst : in std_logic
    );
	
  end component Div_FormConv_Norm;
  
  component Division_pl is
	  generic(
		WN : integer := 16;   --1 integer plus 15 fractional bits
		WD : integer := 16;
		max_shift : integer := 3;  --log2(max(WD,WN))-1  or Width(binary(max(WN,WD))-1
		TWO : integer := 65536;     --2**WN
		PO2WN : integer := 32768;  --2**(WN-1)
		PO2WN2 : integer := 131071  --2**(WN+1)-1
	  );



	  port(
		N_in  : in std_logic_vector(WN-1 downto 0);
		D_in  : in std_logic_vector(WD-1 downto 0);
		sign  : in std_logic;
		bit_shift : in std_logic_vector (max_shift downto 0);
		
		Q_out : out std_logic_vector(WD-1 downto 0):= (others => '0');
		clk : in std_logic;
		rst : in std_logic
	  );
  end component Division_pl; 
  
  
  
begin
  
  UUT1 : Div_FormConv_Norm
    port map (
      N_in     => r_N_in,
      D_in     => r_D_in,
	  sign       => w_sign,
	  bit_shift  => w_bit_shift,
	  N_out    => w_N_out,
	  D_out    => w_D_out,
      clk      => r_clk,
	  rst      => r_rst
      );
   
   UUT2 : Division_pl
    port map (
      rst     => r_rst,
	  clk     => r_clk,
	  N_in    => w_N_out,
	  D_in    => w_D_out,
	  sign    => w_sign,
	  bit_shift => w_bit_shift,
	  Q_out   => w_Q_out
      );
 
  p_clk_gen : process is
    begin 
	  wait for c_clk_period/2;
	  r_clk <= not(r_clk);
  end process p_clk_gen;
	
	
  
	
  process
  FILE file_out : TEXT IS OUT "dataout.txt";
  VARIABLE line_out : LINE;
  VARIABLE output_tmp : INTEGER;
  begin
	
	    r_N_in <= "0110000100000011";
    r_D_in <= "0111000101010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000111010101010";
    r_D_in <= "1010011110010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111110011110";
    r_D_in <= "0111101001100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110001110011";
    r_D_in <= "1000100111001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011101011010";
    r_D_in <= "0101100000100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111001011000000";
    r_D_in <= "0101101100111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111111000011";
    r_D_in <= "0100000000111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100011010011100";
    r_D_in <= "0110111110011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001011111011";
    r_D_in <= "0110110111111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001100100010";
    r_D_in <= "1000000011101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101100111101011";
    r_D_in <= "0111011010010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011111000100";
    r_D_in <= "0100100001110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011100100101110";
    r_D_in <= "1000101000100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110111110010";
    r_D_in <= "1000001001101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100100001110110";
    r_D_in <= "0110000100101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000100101100";
    r_D_in <= "0111000000000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101101000010";
    r_D_in <= "1000010001011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101101110000";
    r_D_in <= "0010100011101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001001001111";
    r_D_in <= "1001011011011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111110101000";
    r_D_in <= "0101010000100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100111111000";
    r_D_in <= "0101000000101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011011011011";
    r_D_in <= "0100101001000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011001000110";
    r_D_in <= "1010001010011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101001000011";
    r_D_in <= "0101000100001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001000000001";
    r_D_in <= "1000111101110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100100001110";
    r_D_in <= "0101100000110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000100110110000";
    r_D_in <= "0110011000011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101010011011";
    r_D_in <= "1010000101111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000000000100100";
    r_D_in <= "1010101110000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100010100100";
    r_D_in <= "0111000010001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110001101101010";
    r_D_in <= "0110010001111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100100100111";
    r_D_in <= "0111110110100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000000110111";
    r_D_in <= "0111010111000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110001101111001";
    r_D_in <= "0110001011010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110101110101";
    r_D_in <= "0011111111001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011100010100100";
    r_D_in <= "0011100110111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101000110100";
    r_D_in <= "0111111000010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000111100001";
    r_D_in <= "0111100110111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000001010101";
    r_D_in <= "0111011000011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011011000001";
    r_D_in <= "0010111001111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100001110111";
    r_D_in <= "0110010011000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100000111011100";
    r_D_in <= "1000110111110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000000001110";
    r_D_in <= "0101001101111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110101101111100";
    r_D_in <= "0110111000111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010110000100";
    r_D_in <= "0101110011011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100101000000";
    r_D_in <= "0010100110110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110000101000100";
    r_D_in <= "0110001101101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001100100011011";
    r_D_in <= "0001101111000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000111111001011";
    r_D_in <= "0111000011001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001011111011";
    r_D_in <= "0111110111011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001110001001";
    r_D_in <= "1001000001010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010011011110";
    r_D_in <= "0110000111110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011110110001";
    r_D_in <= "0111001111101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110011101001";
    r_D_in <= "0001110110001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100100000100";
    r_D_in <= "0011101100010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011101011010";
    r_D_in <= "0110110000000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011111111100";
    r_D_in <= "0111110000110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001101101100100";
    r_D_in <= "1001101110010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110001111010";
    r_D_in <= "0100110011101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111000010101";
    r_D_in <= "0011010010100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100001100001";
    r_D_in <= "1000101100001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001001100111";
    r_D_in <= "1001001000101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111110000001";
    r_D_in <= "0111101000000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010011110110111";
    r_D_in <= "1000000001010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000110000111";
    r_D_in <= "0011000111001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011100110010";
    r_D_in <= "0111111010100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111000001110";
    r_D_in <= "1000110110111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000011010101";
    r_D_in <= "0010000101011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000100111011";
    r_D_in <= "0100000110001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101100101111101";
    r_D_in <= "1000101111101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110001011111110";
    r_D_in <= "0001111001010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101010110110000";
    r_D_in <= "0011010010110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111011101010";
    r_D_in <= "0111001110001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100110101001";
    r_D_in <= "0111101100011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110101000110101";
    r_D_in <= "1000001011011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000010010110";
    r_D_in <= "0110100011001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100011000100";
    r_D_in <= "0010100011000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010111001000";
    r_D_in <= "1010001000011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011000011101";
    r_D_in <= "0100100001100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001110100101";
    r_D_in <= "0110110101111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011111000110";
    r_D_in <= "0010111101010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111001010001";
    r_D_in <= "0111000010101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110100101001100";
    r_D_in <= "0110101010011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011100010000";
    r_D_in <= "0100011001111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111110110100100";
    r_D_in <= "0101111011110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001001011101";
    r_D_in <= "0111001111011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010111010101";
    r_D_in <= "0101111100010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110000101000";
    r_D_in <= "0111000010110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010111011011";
    r_D_in <= "0110010101111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010100001100";
    r_D_in <= "0110110011011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000100010110001";
    r_D_in <= "0110001001111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111010101001";
    r_D_in <= "1000000010000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010000100111";
    r_D_in <= "1010101101100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110010100110";
    r_D_in <= "0100111101000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000011101010";
    r_D_in <= "0101000111000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111100110011";
    r_D_in <= "0101110100100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100101011011";
    r_D_in <= "0001001010101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110010011101";
    r_D_in <= "0010000000011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101100001111";
    r_D_in <= "0110100000001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010010001101";
    r_D_in <= "0101111100111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010110001010";
    r_D_in <= "0101110010100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110110001011001";
    r_D_in <= "0011001011110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010010110100";
    r_D_in <= "0011110110100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100100111011010";
    r_D_in <= "0110010001010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001101000010";
    r_D_in <= "0111001001000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001111011000";
    r_D_in <= "0111111001110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011011111011";
    r_D_in <= "0101110110000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100001011001";
    r_D_in <= "0110100010101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000000101111100";
    r_D_in <= "1010011001111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011100100010";
    r_D_in <= "0110011100100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010000110001";
    r_D_in <= "1001001011110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010010111111";
    r_D_in <= "0100110101110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010001111000";
    r_D_in <= "0111111001110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000111110000";
    r_D_in <= "0101001111111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100111101000";
    r_D_in <= "0110000010111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111111101011";
    r_D_in <= "0001110010110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111101110100";
    r_D_in <= "0110100111000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000010101101";
    r_D_in <= "0001010100111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110011100001";
    r_D_in <= "1000110000001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010010001100";
    r_D_in <= "1001111110001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101000110101";
    r_D_in <= "0101110111101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001011110001010";
    r_D_in <= "1001111011100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001111000111";
    r_D_in <= "0111010000010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011001000111";
    r_D_in <= "0110101111000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001011011000";
    r_D_in <= "1010100000000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101110010100";
    r_D_in <= "0111110110001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010010110111";
    r_D_in <= "0110111001001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100011011010";
    r_D_in <= "0001100111110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110101011111";
    r_D_in <= "0101101101101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011010010100";
    r_D_in <= "0101101010100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010101110110";
    r_D_in <= "1001011111010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111011101111";
    r_D_in <= "1001011000011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011100011010";
    r_D_in <= "1000000011010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000100011101";
    r_D_in <= "0011010111001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010011110111";
    r_D_in <= "0111001100110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111111000111";
    r_D_in <= "0101000010001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001110011010";
    r_D_in <= "0010110100101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001100100001000";
    r_D_in <= "0111111101110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101010111100";
    r_D_in <= "0001010010111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000011001111";
    r_D_in <= "0111010001111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010001100110";
    r_D_in <= "1000000010011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000110111101000";
    r_D_in <= "0111001100001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101101101111";
    r_D_in <= "0111110110101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111100011000";
    r_D_in <= "1001001001000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101000010000";
    r_D_in <= "1000111001011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010010101110";
    r_D_in <= "1000100000001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111011100111";
    r_D_in <= "0110001000110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010111111100";
    r_D_in <= "0100101000001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001111010000000";
    r_D_in <= "0110000111110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010111000000";
    r_D_in <= "0111101011011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101100100001110";
    r_D_in <= "0101111001011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010011000110";
    r_D_in <= "0111100000010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101011001101";
    r_D_in <= "0101011101110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000001000111";
    r_D_in <= "0011010111100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000000000000100";
    r_D_in <= "0100100111000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100111110000";
    r_D_in <= "0111011000011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100001000101";
    r_D_in <= "0010101101011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010011011110";
    r_D_in <= "0101110110010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000011101001";
    r_D_in <= "0011100110110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110100111001";
    r_D_in <= "0111010010000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010001110110";
    r_D_in <= "0101001010000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010111111101";
    r_D_in <= "0110100001001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010111010101";
    r_D_in <= "0111011100000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000100011111";
    r_D_in <= "0101010001110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001100111110110";
    r_D_in <= "0101100001001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101001001101";
    r_D_in <= "0101000011111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111011000101";
    r_D_in <= "0101001111110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010011100101";
    r_D_in <= "0101011101101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110001100010";
    r_D_in <= "1001010111111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100000100100";
    r_D_in <= "0001100101110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110111101100";
    r_D_in <= "0100001100110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011001101100";
    r_D_in <= "0101111100110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011000010101";
    r_D_in <= "0111111111011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011100111010";
    r_D_in <= "0110110000111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010101100011";
    r_D_in <= "0100001011110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101100000011";
    r_D_in <= "0111011010110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111110100011";
    r_D_in <= "0101101001101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010101110010";
    r_D_in <= "0011001000100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010110010001";
    r_D_in <= "0010110101010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101010110000011";
    r_D_in <= "0010111000000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111010111101";
    r_D_in <= "0101111101101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000100011010";
    r_D_in <= "0101111010011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111001010001";
    r_D_in <= "0101110111101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101011111011";
    r_D_in <= "0110010001100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110010000001";
    r_D_in <= "1000100011010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101111001000";
    r_D_in <= "0100000110001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000001001000";
    r_D_in <= "0110010100001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001001010001";
    r_D_in <= "0101000100000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100110100001";
    r_D_in <= "0100100110110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011100010010111";
    r_D_in <= "0111110001000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001110110011";
    r_D_in <= "1000110011110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111100001100";
    r_D_in <= "1001001000010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101001111110";
    r_D_in <= "0100110111101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100001110101";
    r_D_in <= "0100111011110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001100101111";
    r_D_in <= "0100011110110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011011100011";
    r_D_in <= "0111110110001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101000111010";
    r_D_in <= "1001001010010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010010001101";
    r_D_in <= "0101011110111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111100110101";
    r_D_in <= "0000100001100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011001110110";
    r_D_in <= "0101111011011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100001111100";
    r_D_in <= "0101010101011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001001001100100";
    r_D_in <= "0101100000011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100000001011";
    r_D_in <= "0110101101010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000010100010";
    r_D_in <= "0101011110010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111111010001";
    r_D_in <= "0100000101001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110111110001";
    r_D_in <= "1001011101001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111100001011";
    r_D_in <= "0110000110100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010111111001";
    r_D_in <= "0111111011001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001011010010101";
    r_D_in <= "0111100010000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101000110011";
    r_D_in <= "0110011100111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011001000001";
    r_D_in <= "0100011111011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110110101011110";
    r_D_in <= "0010101001010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101110010111";
    r_D_in <= "0011011010101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111110101000001";
    r_D_in <= "0101111101110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110101101001110";
    r_D_in <= "1000101001010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110000110100";
    r_D_in <= "0101001010000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010101011100";
    r_D_in <= "0111101111000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000101110011";
    r_D_in <= "0101000010100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110001101101";
    r_D_in <= "1000010001101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111111100010";
    r_D_in <= "1000111101011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011000111101";
    r_D_in <= "1001110001010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010101001111";
    r_D_in <= "1001011010011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001110000001";
    r_D_in <= "1010011010001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011111110011";
    r_D_in <= "0110100100101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100001001001";
    r_D_in <= "1000110111111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111100011011";
    r_D_in <= "0010111101011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000110100001110";
    r_D_in <= "0100010100111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011000001110";
    r_D_in <= "0101100011111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001011101110";
    r_D_in <= "0101100010110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110101110011001";
    r_D_in <= "1000111011110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101001110101";
    r_D_in <= "0110111101110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110011000000";
    r_D_in <= "1000101000110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100100101110";
    r_D_in <= "1000101000000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101101010011";
    r_D_in <= "0111011001110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100111000010";
    r_D_in <= "0111011101100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101010000100";
    r_D_in <= "1001000100010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010110110100";
    r_D_in <= "0100110101111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100110001010";
    r_D_in <= "0110000110111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010000011010";
    r_D_in <= "1001011001111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110001111000";
    r_D_in <= "0101010101011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101110100110100";
    r_D_in <= "0110011101110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111001101111";
    r_D_in <= "0101101010011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010010001011";
    r_D_in <= "0111011010111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000000101111100";
    r_D_in <= "0011010001110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001000101110";
    r_D_in <= "0111110111000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101111010111";
    r_D_in <= "0110110011010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110001001000";
    r_D_in <= "0101010001011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001110000010";
    r_D_in <= "0110000110011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101100100001011";
    r_D_in <= "1000110011101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000111101101000";
    r_D_in <= "1000010111100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000110001001010";
    r_D_in <= "0111111101101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000100101001001";
    r_D_in <= "0101100111101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111001011010101";
    r_D_in <= "0101011111001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010000100011";
    r_D_in <= "1000001001101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010110011110";
    r_D_in <= "1000000111100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010111101101";
    r_D_in <= "1000010101111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111101101010";
    r_D_in <= "0110100000101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011110110101";
    r_D_in <= "0100110100000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111011000001";
    r_D_in <= "0110101100001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101100011011110";
    r_D_in <= "0110001010011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000100001000";
    r_D_in <= "0011001101010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101110000101";
    r_D_in <= "0100100011101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101110101101000";
    r_D_in <= "0100010001001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000110001100011";
    r_D_in <= "1000011100001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110101111010101";
    r_D_in <= "0101000001000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010101100111";
    r_D_in <= "1000101000001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010011000111";
    r_D_in <= "0110000111001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000010010010";
    r_D_in <= "0101000010011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101101110010";
    r_D_in <= "0001111010110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111010000001";
    r_D_in <= "0101101001111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111011001111";
    r_D_in <= "0110111011111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111011111110";
    r_D_in <= "0010000011011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100010101110";
    r_D_in <= "0110100010110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010010000000";
    r_D_in <= "1000100100011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011111000000";
    r_D_in <= "0101101000110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110001011101";
    r_D_in <= "1000011101000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001011011100";
    r_D_in <= "1010111110100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110111010011";
    r_D_in <= "0011000011111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111111110010";
    r_D_in <= "0101111010001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111100110101";
    r_D_in <= "1000010111110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011110010010";
    r_D_in <= "0111010010100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001000110010";
    r_D_in <= "0111111101101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110001010110";
    r_D_in <= "0111001001000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010100100111";
    r_D_in <= "0111011010011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011100001001";
    r_D_in <= "0110100101001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011001000111";
    r_D_in <= "0110110010010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111010010011";
    r_D_in <= "0111110110100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111111110000";
    r_D_in <= "0110011000011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000010011110";
    r_D_in <= "0101111000111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010010000010";
    r_D_in <= "0010001100101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010001111100";
    r_D_in <= "0011101110100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100101000000";
    r_D_in <= "0111111001001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011101111011";
    r_D_in <= "1001101011010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000110100111";
    r_D_in <= "0101001001110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111110010100";
    r_D_in <= "1000110001001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011011111011";
    r_D_in <= "0100011110110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111001110101010";
    r_D_in <= "0100110000101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111010001100";
    r_D_in <= "0111010110101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001000100111";
    r_D_in <= "0011111101010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001000100001";
    r_D_in <= "0111101110101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110001000100";
    r_D_in <= "0100110010010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011011011110";
    r_D_in <= "0101011011110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010010010001";
    r_D_in <= "0101010001110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001001111000";
    r_D_in <= "0001100100000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111100111011";
    r_D_in <= "0101011101001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010111100111";
    r_D_in <= "0110001101101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011111111011";
    r_D_in <= "0101100011111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001000000001001";
    r_D_in <= "0111011100101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001010001101110";
    r_D_in <= "0110111111011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101101111011";
    r_D_in <= "0111001100000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111100001101";
    r_D_in <= "0110100011110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011100101001";
    r_D_in <= "1000101101001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001111000111111";
    r_D_in <= "0110000111110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100011111011101";
    r_D_in <= "0011101110111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111011100000";
    r_D_in <= "0001000111010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100000000100";
    r_D_in <= "1000010011100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101101000001";
    r_D_in <= "0010000110011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001101100100";
    r_D_in <= "1001111101100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001100000101";
    r_D_in <= "0110010001101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010001010001010";
    r_D_in <= "0111111101111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101101010011";
    r_D_in <= "0010100000001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110001110111110";
    r_D_in <= "0110010110000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110100111100";
    r_D_in <= "0111111010011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111011011000";
    r_D_in <= "0111111011110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010110110110";
    r_D_in <= "0101101001011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101001101000";
    r_D_in <= "0100101001101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111000101110";
    r_D_in <= "1001000011001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101001100011";
    r_D_in <= "0100101110101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011111001100";
    r_D_in <= "1001000111111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111001100011";
    r_D_in <= "0111011011001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110111111101";
    r_D_in <= "0100001000111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011111110100";
    r_D_in <= "0100110110111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001100111000";
    r_D_in <= "0101001100111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100010110010";
    r_D_in <= "1001100101011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101100010011";
    r_D_in <= "0011111000100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100110110010";
    r_D_in <= "0111111010101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100011110011";
    r_D_in <= "0010100110001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001001010000";
    r_D_in <= "1001010000100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101110100100";
    r_D_in <= "0111011101011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000110010000110";
    r_D_in <= "0001111100011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000111000000";
    r_D_in <= "0011010101001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000000100101";
    r_D_in <= "0110110101001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000110101001010";
    r_D_in <= "0111111100100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111001001111110";
    r_D_in <= "0111100001110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110110100110";
    r_D_in <= "0111001011100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111000011110";
    r_D_in <= "0010011011001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011010110001";
    r_D_in <= "0101011111100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011001110101";
    r_D_in <= "1001010001000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011011110110011";
    r_D_in <= "0011011111011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010010001111";
    r_D_in <= "0111110110001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001011011101111";
    r_D_in <= "0100010001011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100101010001";
    r_D_in <= "0100100100010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111000111101011";
    r_D_in <= "1010101100111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001000011111";
    r_D_in <= "0100100011010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011010000010";
    r_D_in <= "1000011011011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110101001100";
    r_D_in <= "0111000111110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011100000111011";
    r_D_in <= "0100101001100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011000001101";
    r_D_in <= "0001111011001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111100110001";
    r_D_in <= "0101001111001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100110101010";
    r_D_in <= "0101000011100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100100001001001";
    r_D_in <= "0100101010010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000000011000111";
    r_D_in <= "1000011101110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101010011110";
    r_D_in <= "0101111100111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110101110000111";
    r_D_in <= "0011101101010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100010000111";
    r_D_in <= "0101100001101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110001011011";
    r_D_in <= "1001000011111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010100011111";
    r_D_in <= "1000000110001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011011101000";
    r_D_in <= "0100110000000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110010000111";
    r_D_in <= "0010110111010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111000001000";
    r_D_in <= "0110001110101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110101110011";
    r_D_in <= "0111100000101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101000001001";
    r_D_in <= "1000010000110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110010010101";
    r_D_in <= "0100001000101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111100101111";
    r_D_in <= "0110001000010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000000000101111";
    r_D_in <= "1000010101101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111100101011";
    r_D_in <= "0100100110000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010011001110";
    r_D_in <= "1001111011011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111111011111";
    r_D_in <= "0101000000100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101010010111";
    r_D_in <= "1010100000111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010101011101";
    r_D_in <= "0100111101111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010011101100";
    r_D_in <= "0111010011110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100011101010000";
    r_D_in <= "1000101101001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111011011111";
    r_D_in <= "0110011011000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100011111000";
    r_D_in <= "0101111111001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101010110100";
    r_D_in <= "0000101010111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110111100110";
    r_D_in <= "0010000100010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010001110011";
    r_D_in <= "0011010000010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000111000010";
    r_D_in <= "1001011001101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011100000011";
    r_D_in <= "0010101100111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001000011110111";
    r_D_in <= "1001111111100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101101001011";
    r_D_in <= "0010111111001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100011001001111";
    r_D_in <= "0111011011110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100011110101011";
    r_D_in <= "1000001010111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001000110101011";
    r_D_in <= "1000111000011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100100110010";
    r_D_in <= "0111011101001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111011100110";
    r_D_in <= "0011011100110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000011001100";
    r_D_in <= "0101011001011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000000011111";
    r_D_in <= "0110101101001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011010001101";
    r_D_in <= "0010110111001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011011011000000";
    r_D_in <= "0011011110011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100110111011110";
    r_D_in <= "0110001001110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111100010100";
    r_D_in <= "0011111111001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101100001101";
    r_D_in <= "0001101011101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101101101100";
    r_D_in <= "1010101101011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001101000010";
    r_D_in <= "1010100111010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000011010111";
    r_D_in <= "0110101110000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000000000101";
    r_D_in <= "0001000001001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001111011011";
    r_D_in <= "0111111001000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101100101000";
    r_D_in <= "0100000110010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000010101011";
    r_D_in <= "0011100110011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000010000010";
    r_D_in <= "0110100001111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011110101100";
    r_D_in <= "0101001010010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001000000101";
    r_D_in <= "0100111001110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010100000000";
    r_D_in <= "0011011000000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000110101000";
    r_D_in <= "0101011001111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110000111010";
    r_D_in <= "0110010000010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001111000010";
    r_D_in <= "1001011000010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010110011101";
    r_D_in <= "0111100100101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010010110110";
    r_D_in <= "1010100000101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111110100110";
    r_D_in <= "0111011111101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010100010001";
    r_D_in <= "0101110001010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001001111111111";
    r_D_in <= "0100100100010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110111010100";
    r_D_in <= "1000111000110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101111111000";
    r_D_in <= "1001000000001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000001100100";
    r_D_in <= "0111010011000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010001100010010";
    r_D_in <= "0011000100101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101100111000";
    r_D_in <= "0111100010111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100001111001";
    r_D_in <= "0010100010000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100111110110";
    r_D_in <= "0110011000011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101001000001";
    r_D_in <= "0110010001010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000011111101";
    r_D_in <= "0110100110111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100010101110";
    r_D_in <= "0011011010111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110101111011001";
    r_D_in <= "1000000011010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010010111001";
    r_D_in <= "0100001001000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011101000100";
    r_D_in <= "0100011101011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111100010100";
    r_D_in <= "0101010010011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010111010011";
    r_D_in <= "0111111011011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101110100001";
    r_D_in <= "0100110000100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110101100010";
    r_D_in <= "1011000110011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101000001000000";
    r_D_in <= "0011101001101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000111111101";
    r_D_in <= "0110010011001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011101101001";
    r_D_in <= "0110001011000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011100100101010";
    r_D_in <= "0100011000111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110010001101";
    r_D_in <= "0110000111101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111001011100";
    r_D_in <= "0110011110000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010011010111110";
    r_D_in <= "0110011111010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011000111101";
    r_D_in <= "0110101110000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101101000111";
    r_D_in <= "1001100011001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001111011011";
    r_D_in <= "0110111001100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011111100001";
    r_D_in <= "0111100100001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110011111000";
    r_D_in <= "0111001010110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010010101001";
    r_D_in <= "0111110100110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110000111001";
    r_D_in <= "0111001010001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001011000110011";
    r_D_in <= "1001000101010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001111000111000";
    r_D_in <= "0111000000000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101100010010";
    r_D_in <= "1000011011100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101001101011";
    r_D_in <= "0101001111011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100001111000";
    r_D_in <= "0010111100000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011100100010";
    r_D_in <= "0101101011011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111010010000";
    r_D_in <= "1000010110101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100011100101";
    r_D_in <= "1010000001100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010100101010";
    r_D_in <= "1001010101011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110110001101000";
    r_D_in <= "0001001111000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101000000101000";
    r_D_in <= "0101000101011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110001110110110";
    r_D_in <= "1001110100001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111101110111";
    r_D_in <= "0010001001010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001011100101110";
    r_D_in <= "0011100100110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110100000111111";
    r_D_in <= "0110100001010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001001110000";
    r_D_in <= "0110111100100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001011101100010";
    r_D_in <= "1000101010011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010001100000011";
    r_D_in <= "1000000100101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000111011001";
    r_D_in <= "0110110111010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110101110000001";
    r_D_in <= "0110101110101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111110111101";
    r_D_in <= "1001101101000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010110001011";
    r_D_in <= "0111010100111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000111111111111";
    r_D_in <= "0111000010001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010010110110";
    r_D_in <= "0110001100100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110011100011";
    r_D_in <= "0101010110000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000010111110";
    r_D_in <= "0010101011101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011011110100001";
    r_D_in <= "0011100110000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111000010111";
    r_D_in <= "0111101001110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011111011110";
    r_D_in <= "0010011101011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011001110111";
    r_D_in <= "0011001011010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010101000110011";
    r_D_in <= "0010110000010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101111000010";
    r_D_in <= "0011111110110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011000100101";
    r_D_in <= "0111110111011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010100110111";
    r_D_in <= "0111100000101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000001111101";
    r_D_in <= "1000100111001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110101111110110";
    r_D_in <= "0010010011100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110101001101110";
    r_D_in <= "1010010001111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001101100001";
    r_D_in <= "0100000100011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001010001100";
    r_D_in <= "0000111100000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000010001110";
    r_D_in <= "0011100010001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111110110010";
    r_D_in <= "1000011010010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100010000100";
    r_D_in <= "0101101000111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101100111001";
    r_D_in <= "0110011010000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111100001000";
    r_D_in <= "0011001010110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010001100001";
    r_D_in <= "1000011101101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101000000101";
    r_D_in <= "0111111110011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111010100110";
    r_D_in <= "0100000101100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000011010011";
    r_D_in <= "1000100011111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001011110001011";
    r_D_in <= "0110101000110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001110001011";
    r_D_in <= "0100000011001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001101001111";
    r_D_in <= "1000000011111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010010000101";
    r_D_in <= "0010101111100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110001100110";
    r_D_in <= "1001000000100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001111001001";
    r_D_in <= "0100010001011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001001010000";
    r_D_in <= "0100001011001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101110000110";
    r_D_in <= "0110011000001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100011010010";
    r_D_in <= "0111111111001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001101001000110";
    r_D_in <= "0110100011110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001001001000";
    r_D_in <= "0111000110011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100000010000110";
    r_D_in <= "0100010000100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011001000000";
    r_D_in <= "0111100011100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100001101010000";
    r_D_in <= "0101110101000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001100111001011";
    r_D_in <= "0001110000001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111111100101";
    r_D_in <= "0101001110011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110010000001";
    r_D_in <= "0110110001111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000111110100";
    r_D_in <= "0100110110010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001100000111101";
    r_D_in <= "0011001000101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001100010001";
    r_D_in <= "0000010000110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011011110100";
    r_D_in <= "0110100100101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010011011100";
    r_D_in <= "0101000001000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000110010011";
    r_D_in <= "0101010100100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111110001110100";
    r_D_in <= "0000010001011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110101000011000";
    r_D_in <= "0110110000010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010100000000";
    r_D_in <= "0111010111000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101010010111";
    r_D_in <= "0101000001100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000110101001";
    r_D_in <= "0110010101001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110101101101";
    r_D_in <= "0011001000011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111101100010";
    r_D_in <= "0001001010001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100001000010110";
    r_D_in <= "0101100110011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001111101000";
    r_D_in <= "0101100100110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001010001100";
    r_D_in <= "1000011010110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000001101110";
    r_D_in <= "0111000011001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001011110101111";
    r_D_in <= "0110100001110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100100110111";
    r_D_in <= "1001001001011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101010001001101";
    r_D_in <= "0110001101111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001001001100";
    r_D_in <= "0000001001001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101111111110";
    r_D_in <= "1001000100100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110101000011110";
    r_D_in <= "0001111000011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000101010011";
    r_D_in <= "0011011101100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010000000111";
    r_D_in <= "0110111101000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011011001001";
    r_D_in <= "1000100011010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110001111101011";
    r_D_in <= "0011100111001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000100111001001";
    r_D_in <= "0011001110010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010110011011";
    r_D_in <= "1001000011011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100001111100100";
    r_D_in <= "1000011111011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011001110111";
    r_D_in <= "0000110110000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011010011000";
    r_D_in <= "0000100111101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011100110000";
    r_D_in <= "1000000101110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011011001011";
    r_D_in <= "0010001100000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111001001101";
    r_D_in <= "1000111011000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110111111110";
    r_D_in <= "1001001101010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111100000011";
    r_D_in <= "0100001101010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001010011001";
    r_D_in <= "0100010101010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011110001011";
    r_D_in <= "0100100010000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101011001010";
    r_D_in <= "0100101011101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101010100111";
    r_D_in <= "0010110101111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000110111101100";
    r_D_in <= "0000111001100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100111010110";
    r_D_in <= "1000001011101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110101011111100";
    r_D_in <= "1010001001001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101100001100";
    r_D_in <= "0110011110110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011001000110";
    r_D_in <= "1000110100110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111000001011";
    r_D_in <= "0000111111101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100110010100";
    r_D_in <= "0111001010000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010101011000100";
    r_D_in <= "0111010101010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100101010011";
    r_D_in <= "0001111111011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011101101101";
    r_D_in <= "0100000001111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101110000001";
    r_D_in <= "0110100100010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111100110111";
    r_D_in <= "0001011100101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100111000010";
    r_D_in <= "0111100100101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010000011100";
    r_D_in <= "0111000010101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101110110110";
    r_D_in <= "0100001000101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011010101111";
    r_D_in <= "0111110101001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110111101110";
    r_D_in <= "1001011110110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000100000001";
    r_D_in <= "0110001110110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010100000101";
    r_D_in <= "1010010101101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010011101111";
    r_D_in <= "1010000100100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001011001011";
    r_D_in <= "0101111100110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101000010010";
    r_D_in <= "0010001101110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000110010001011";
    r_D_in <= "0011000000011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101010011111";
    r_D_in <= "0100000100110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100101100011";
    r_D_in <= "0110001001110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000101001101";
    r_D_in <= "0100111001110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000111111011";
    r_D_in <= "0101110100111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110001101011001";
    r_D_in <= "0111001101001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111010000011";
    r_D_in <= "0011000100101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001111001001";
    r_D_in <= "0101111001001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101110000000";
    r_D_in <= "0100111111011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000101100000";
    r_D_in <= "0111000100011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110000100111";
    r_D_in <= "1000011001111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011100010101";
    r_D_in <= "1010101101100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010101101010";
    r_D_in <= "0110001111100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110001000010";
    r_D_in <= "0110111000100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010101011000";
    r_D_in <= "0111101010111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110010001000";
    r_D_in <= "1011001001110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010111000101";
    r_D_in <= "0111010101010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101000001111";
    r_D_in <= "0111101000010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111001011011";
    r_D_in <= "0110111010011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101011111100";
    r_D_in <= "0011100100110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111011100101";
    r_D_in <= "0111010101100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100111000100";
    r_D_in <= "0110111101000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010110001111";
    r_D_in <= "0110010111110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110000100010111";
    r_D_in <= "0110001010010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010001111001110";
    r_D_in <= "1001010000011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100101101000";
    r_D_in <= "0111011111101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100011111000";
    r_D_in <= "0100100110010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110110101001";
    r_D_in <= "0101011100110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001011101011";
    r_D_in <= "1000110000111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010101011001";
    r_D_in <= "0000100010100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100100100011";
    r_D_in <= "0010111110101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111111111101";
    r_D_in <= "0111111001100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101001010001";
    r_D_in <= "1001010111000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100000010110";
    r_D_in <= "0111101010111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011100100010";
    r_D_in <= "1010000101100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101100111100";
    r_D_in <= "0010010011110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011101110011";
    r_D_in <= "0111101100000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001110101000";
    r_D_in <= "0110111000101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011000001001011";
    r_D_in <= "1001010101010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011101111011";
    r_D_in <= "0110011000110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101001011011";
    r_D_in <= "0010111011110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001011010000101";
    r_D_in <= "0110111001010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110110100101";
    r_D_in <= "0110110110101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000100110100";
    r_D_in <= "0101111111011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100000000111";
    r_D_in <= "1000110101101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110101000100";
    r_D_in <= "0101001110100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010010110011";
    r_D_in <= "0110001010011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011011000010111";
    r_D_in <= "0011011101000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111111010001";
    r_D_in <= "0101000110100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110100010000110";
    r_D_in <= "0111111010101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010001010010001";
    r_D_in <= "0111001011100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010101101000";
    r_D_in <= "1001001100101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001111111111101";
    r_D_in <= "0110000011111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111000001111";
    r_D_in <= "1010100001110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100110010010111";
    r_D_in <= "0101111010110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010101011011";
    r_D_in <= "0101110100001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000000000110";
    r_D_in <= "0100011010011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000011001011";
    r_D_in <= "0110000111100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010010011110";
    r_D_in <= "0110110101111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001111000111";
    r_D_in <= "0011001111010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011010010000";
    r_D_in <= "0101000110001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010110101001";
    r_D_in <= "0001011011000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000111011011101";
    r_D_in <= "1000101111111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100001001110";
    r_D_in <= "0111110001110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010100100111";
    r_D_in <= "1000111111111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111100001111";
    r_D_in <= "1001111010011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100101010010";
    r_D_in <= "0110010101010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100011111001";
    r_D_in <= "0011001001000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101001111010";
    r_D_in <= "0100110100110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111111011110";
    r_D_in <= "0111110100110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100000011101010";
    r_D_in <= "1000001100010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100010001110";
    r_D_in <= "0011110110110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000110011001";
    r_D_in <= "0110110010001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100011011100";
    r_D_in <= "1000001100111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001011111010110";
    r_D_in <= "1001101000011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000101011101";
    r_D_in <= "1001011111000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001010000011";
    r_D_in <= "0100001010010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010100000010";
    r_D_in <= "0111100111000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111110101101";
    r_D_in <= "0111111010100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111111110000";
    r_D_in <= "0111100011100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101000111000000";
    r_D_in <= "0100001001101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001101010111";
    r_D_in <= "1000010001001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100101110110";
    r_D_in <= "0101111001001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100111100100";
    r_D_in <= "1000111001011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010001000101100";
    r_D_in <= "0011111011110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111001001001010";
    r_D_in <= "0011000000011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111100011110";
    r_D_in <= "0111110001101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011011001010101";
    r_D_in <= "1000010010011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110100011000";
    r_D_in <= "0110110100110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011111011100";
    r_D_in <= "1000111111011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000110000111";
    r_D_in <= "0010001101001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000000011100";
    r_D_in <= "0101010110000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011010100010";
    r_D_in <= "0011111010000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100000100110110";
    r_D_in <= "0110101011111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111001010110111";
    r_D_in <= "0011011001110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100011110011";
    r_D_in <= "0011111010111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110110010100011";
    r_D_in <= "0011110011000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110010001000";
    r_D_in <= "0010111010111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101110101110";
    r_D_in <= "1001101011011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000111010001100";
    r_D_in <= "0111001000101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111111011100";
    r_D_in <= "1010010011100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100010001000";
    r_D_in <= "0101100111110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011101011000";
    r_D_in <= "0000111010001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110100111011";
    r_D_in <= "0101011011010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010100100000";
    r_D_in <= "0011000011011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100001000010110";
    r_D_in <= "1000101111011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010101010001";
    r_D_in <= "1010101111111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100001001100";
    r_D_in <= "0111001000101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111001111000";
    r_D_in <= "0001001101001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011101111100";
    r_D_in <= "0100111100110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010101100000";
    r_D_in <= "0010001010000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110011001111";
    r_D_in <= "0101100111110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100101101101";
    r_D_in <= "0011111000101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001000001010";
    r_D_in <= "0011100110000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100000110110010";
    r_D_in <= "0100000111001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111011010110";
    r_D_in <= "1000000011110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011010011011";
    r_D_in <= "0010100110010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101111001000";
    r_D_in <= "0111111010011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000110011010010";
    r_D_in <= "1000010101010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010111101111";
    r_D_in <= "1000000000011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110110110011";
    r_D_in <= "0100100100101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110000111100";
    r_D_in <= "0001110101110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000101001110";
    r_D_in <= "0110001101100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001000000101111";
    r_D_in <= "0111001110100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111000000001000";
    r_D_in <= "0111110010011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011011011010010";
    r_D_in <= "0100001101100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110001101111010";
    r_D_in <= "0110101010011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100011101010";
    r_D_in <= "0111101110100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011111011101";
    r_D_in <= "1000101001110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110011110101";
    r_D_in <= "1000001101101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101011000010";
    r_D_in <= "0101110111101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011101101011";
    r_D_in <= "0111101100011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010111010010";
    r_D_in <= "0100101100110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010001111111";
    r_D_in <= "0111111110001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101101001000";
    r_D_in <= "0101100100101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111110010010";
    r_D_in <= "0110001101011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111110111101";
    r_D_in <= "1000110011010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110110100010000";
    r_D_in <= "0111000110010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011011010100";
    r_D_in <= "0011000110001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010000101111";
    r_D_in <= "0011101100110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101011100001";
    r_D_in <= "0011111111000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011100000001000";
    r_D_in <= "0111011100001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011001101111";
    r_D_in <= "0101000111100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010001100101100";
    r_D_in <= "0111100110001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110101001010";
    r_D_in <= "0110010010100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001000111011";
    r_D_in <= "0110000010001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101101001000";
    r_D_in <= "0110111001110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010010101000";
    r_D_in <= "0111001001010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110001110111001";
    r_D_in <= "0010110101101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000110100000101";
    r_D_in <= "0110000101100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000101000110";
    r_D_in <= "0101110100000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110001110100010";
    r_D_in <= "1000001011110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111010100110";
    r_D_in <= "0111111001100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110001010101";
    r_D_in <= "0111000100101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110100000110101";
    r_D_in <= "1001111111010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000001111010";
    r_D_in <= "0010011011010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011000001011";
    r_D_in <= "1000100010010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101101101110";
    r_D_in <= "0011110001010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010000101100";
    r_D_in <= "1000101011000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001000011101011";
    r_D_in <= "1001100101101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101110011010011";
    r_D_in <= "0111111011111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101110010011001";
    r_D_in <= "0101110110001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000111101001";
    r_D_in <= "0111000101110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111001011000010";
    r_D_in <= "0101100011011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001000001100011";
    r_D_in <= "1010001101011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010011011011";
    r_D_in <= "0101110110010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111011101011";
    r_D_in <= "1001110111000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011001001000";
    r_D_in <= "0100001001001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010000111011";
    r_D_in <= "1001110011011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101100010101";
    r_D_in <= "0111010000001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001100011000000";
    r_D_in <= "0110110010100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110100101010011";
    r_D_in <= "1001111101100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100001010111";
    r_D_in <= "0111100001101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010110101010";
    r_D_in <= "0101001010011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101110101111";
    r_D_in <= "0101110011000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111011111001";
    r_D_in <= "1000111000110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110000110011";
    r_D_in <= "0110110100011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111001111011";
    r_D_in <= "0110101100010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111001010101";
    r_D_in <= "0101111011011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001011101110";
    r_D_in <= "0101011100101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101101110000";
    r_D_in <= "0111001001001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111000111000001";
    r_D_in <= "1000010011101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000000100011";
    r_D_in <= "0101111001000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101111011000";
    r_D_in <= "1000010101001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011110110111";
    r_D_in <= "0101110001001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100111000010";
    r_D_in <= "0111011000011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111000101000";
    r_D_in <= "1010011100101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111101000000";
    r_D_in <= "0001111101001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111100111110";
    r_D_in <= "0101010001011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111001001011";
    r_D_in <= "0110001111001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110010011100";
    r_D_in <= "1000101001011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101001110101";
    r_D_in <= "0110001001011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000010111000";
    r_D_in <= "1000001100101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101010001100";
    r_D_in <= "0100111100011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001000000101";
    r_D_in <= "0111010000001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001011101011";
    r_D_in <= "0100001111111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100001100000010";
    r_D_in <= "0101010110111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011001001011";
    r_D_in <= "0111001110001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000000110001011";
    r_D_in <= "1000010001011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111111000100";
    r_D_in <= "0110000011001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011101000110";
    r_D_in <= "0111100000111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101101110100";
    r_D_in <= "0101110011100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111110101101";
    r_D_in <= "0011011100111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100011010110";
    r_D_in <= "0110101011111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111010010100";
    r_D_in <= "0011110100001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111000000011";
    r_D_in <= "0011010010111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000001101111";
    r_D_in <= "0010010010010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111000010000";
    r_D_in <= "0101111101111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111111100001";
    r_D_in <= "0011001111111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011101100110";
    r_D_in <= "0111111110001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111110010100";
    r_D_in <= "0111111110001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100000111111010";
    r_D_in <= "0100001110001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000101001010";
    r_D_in <= "0101101001010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101101101101";
    r_D_in <= "0111011000000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010001000111111";
    r_D_in <= "0110111010000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100011110011";
    r_D_in <= "0111100000101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111001001001";
    r_D_in <= "0010100001111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000011000000";
    r_D_in <= "0100011111001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101000111101";
    r_D_in <= "1001100000000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000011100000";
    r_D_in <= "0100010101000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001001011111";
    r_D_in <= "0111010100001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001100010001001";
    r_D_in <= "0001101101111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111011010100";
    r_D_in <= "0101111100000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010110111011";
    r_D_in <= "0110111110101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001101001000";
    r_D_in <= "1000001000101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010110011001";
    r_D_in <= "0100000001111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010100111100";
    r_D_in <= "0111010010101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010110010010";
    r_D_in <= "0001101001110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111010001111";
    r_D_in <= "1000110000110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010001011110";
    r_D_in <= "0111101010001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101010110111";
    r_D_in <= "1001010001001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111111011100";
    r_D_in <= "0111010111011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111010001100";
    r_D_in <= "0010011101000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101111100111";
    r_D_in <= "0110100010101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111000101010";
    r_D_in <= "0111000010111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110101011001";
    r_D_in <= "0111010100011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000110010101100";
    r_D_in <= "0011000010111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001111111011000";
    r_D_in <= "1001100111101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011111101011";
    r_D_in <= "1001000010010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000001111110";
    r_D_in <= "0100001011100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100110011010011";
    r_D_in <= "0100010100010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111100110111";
    r_D_in <= "1000111100111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000110100011010";
    r_D_in <= "1000011011010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010101001100";
    r_D_in <= "0110010111110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000000001101011";
    r_D_in <= "1001110111001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011111000010";
    r_D_in <= "0100111001101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111111000000";
    r_D_in <= "1000011110010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111100111110";
    r_D_in <= "0100110001100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000100100010011";
    r_D_in <= "0001101100000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000001111111";
    r_D_in <= "0110111000101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111000100110";
    r_D_in <= "0110111110000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011110101011";
    r_D_in <= "1000001010101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101110111111";
    r_D_in <= "0111011000011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111010000011";
    r_D_in <= "0110010010100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001011100010101";
    r_D_in <= "0111000011001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010111111011";
    r_D_in <= "0100001100011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001110001101";
    r_D_in <= "0111001110110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101110111010";
    r_D_in <= "1000100010011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000100100011001";
    r_D_in <= "0010110011100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111000100000";
    r_D_in <= "0101111000100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110011000000";
    r_D_in <= "0101110010101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101110001000110";
    r_D_in <= "0110000001111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010011100001";
    r_D_in <= "0110000100010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110000101101100";
    r_D_in <= "0110111110101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011110010110";
    r_D_in <= "0101100111000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100101011000";
    r_D_in <= "0110011101101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110100001111";
    r_D_in <= "0101111010111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110101011100001";
    r_D_in <= "0011101000100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101010111111";
    r_D_in <= "0011000011111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110001110110";
    r_D_in <= "1000010001101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100100010100111";
    r_D_in <= "0110000111000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001111101010";
    r_D_in <= "0110111000011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000111000110";
    r_D_in <= "0111111011010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111110101110";
    r_D_in <= "0110011001101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111110001011";
    r_D_in <= "0111001110000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000100100111";
    r_D_in <= "0010000100110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001101010000001";
    r_D_in <= "1000100011100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001011110111";
    r_D_in <= "0111001010111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010111111101";
    r_D_in <= "0010111011101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111110011101110";
    r_D_in <= "0110010101001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111100101100";
    r_D_in <= "0010011111111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101000111010010";
    r_D_in <= "0010111000110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011001110101";
    r_D_in <= "0010101100110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001101000100";
    r_D_in <= "1000100110100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100111000000";
    r_D_in <= "1010000111001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101000101110";
    r_D_in <= "0011000000010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001110000111";
    r_D_in <= "0011010101110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111001001110";
    r_D_in <= "0110011000111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001011001011100";
    r_D_in <= "0111110101101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100110110110";
    r_D_in <= "1001101000100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010101000100010";
    r_D_in <= "0111000101100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110000110111";
    r_D_in <= "0101110001100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010011010000110";
    r_D_in <= "0100001010100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011101101111";
    r_D_in <= "0101101001011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111010000110";
    r_D_in <= "0000100111001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010111010110";
    r_D_in <= "1000101110010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001001110011";
    r_D_in <= "0110111100001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000110100001110";
    r_D_in <= "0100100100001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111001011110";
    r_D_in <= "0101101011011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001010101000";
    r_D_in <= "0111111010110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101000011000";
    r_D_in <= "0011100100101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010011010000";
    r_D_in <= "1000101110111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100111000110";
    r_D_in <= "0110100100101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011001011010";
    r_D_in <= "0111101100100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101110000000";
    r_D_in <= "0101110110000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111110110100001";
    r_D_in <= "0101100011001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100000010000";
    r_D_in <= "0100010101100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001011010001010";
    r_D_in <= "1000001010000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111101110100";
    r_D_in <= "1000111100110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111011110001";
    r_D_in <= "0111111011111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011001010100";
    r_D_in <= "0011111011000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001011001101001";
    r_D_in <= "0110110011001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011111000000";
    r_D_in <= "1000000100110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101110111000";
    r_D_in <= "1001100011000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000100111101011";
    r_D_in <= "0010101010011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010111011010";
    r_D_in <= "0110011011011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010000011100";
    r_D_in <= "0111111010011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110001111110";
    r_D_in <= "1001010000011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010011011001";
    r_D_in <= "0110101111110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001100010011";
    r_D_in <= "0101011101101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001111000101000";
    r_D_in <= "0111011011101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010011001010";
    r_D_in <= "1000010100001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011011001011";
    r_D_in <= "1001010011101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100100100000001";
    r_D_in <= "0110110000111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101011011000";
    r_D_in <= "1000101010001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010011100100";
    r_D_in <= "1001000110100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000001101101";
    r_D_in <= "0101011000000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100111111111";
    r_D_in <= "0101110111010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110000101111";
    r_D_in <= "0101111011010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011100110111";
    r_D_in <= "0000100011101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101001110101";
    r_D_in <= "0011111101101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110110110010";
    r_D_in <= "0011110111000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111000001101";
    r_D_in <= "0111001101010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001010111101";
    r_D_in <= "0110110101000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001001011101";
    r_D_in <= "0111010011001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111110110010";
    r_D_in <= "0011110111100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001100111000";
    r_D_in <= "0110011000100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001101110001";
    r_D_in <= "0111001000001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111101100111";
    r_D_in <= "0011011011101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111001011100100";
    r_D_in <= "0101001111011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101000111110";
    r_D_in <= "0111110111001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001000101111111";
    r_D_in <= "1000001010000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001010101111";
    r_D_in <= "0100100011011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001111101001100";
    r_D_in <= "0110110000010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000110011101";
    r_D_in <= "0101111011110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011001000001";
    r_D_in <= "0111110101101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110111111110";
    r_D_in <= "0111101011010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010001011001";
    r_D_in <= "0100000111001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111110111010101";
    r_D_in <= "0110001100110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000001001010";
    r_D_in <= "0011111000110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100010010101";
    r_D_in <= "0110100010110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111010110110";
    r_D_in <= "0110101011110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011100000001";
    r_D_in <= "0111010000011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111011101001";
    r_D_in <= "0110011010110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001101001100010";
    r_D_in <= "1001011110001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111110000010";
    r_D_in <= "0001110110010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011010111010";
    r_D_in <= "1000011010101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101000110111";
    r_D_in <= "1000000000011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000110001111";
    r_D_in <= "0110101100101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011001010001";
    r_D_in <= "0000101111011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100100101101";
    r_D_in <= "0110011100110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001000110001";
    r_D_in <= "1000010011101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100111000111";
    r_D_in <= "0111011001010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001011111101";
    r_D_in <= "0110011101110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110001010001";
    r_D_in <= "0111001011101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011000000000000";
    r_D_in <= "0101000101000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000110010110";
    r_D_in <= "0110111110011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101100000100";
    r_D_in <= "1000100110111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110101011001";
    r_D_in <= "0110010101101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011100001110100";
    r_D_in <= "0011100010110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111110100111";
    r_D_in <= "0111111010101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101110011000111";
    r_D_in <= "0011111000011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000010000111";
    r_D_in <= "0110010000110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101100100000";
    r_D_in <= "1000000111111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011010001101";
    r_D_in <= "0010000011100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011001101111";
    r_D_in <= "0110100001000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011011110010111";
    r_D_in <= "0100100011001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101101100011";
    r_D_in <= "0100010101101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001001111010";
    r_D_in <= "0110110110001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101110101011";
    r_D_in <= "0110000011110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101000011011";
    r_D_in <= "0001101101000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011100010010100";
    r_D_in <= "0111101011011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110101110000";
    r_D_in <= "0011010111100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010001100001";
    r_D_in <= "0101010100001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111101011111";
    r_D_in <= "0111101101101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110110111101101";
    r_D_in <= "0111000010001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110110010010101";
    r_D_in <= "0101110111001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001100011111001";
    r_D_in <= "0111111101110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101100100001";
    r_D_in <= "0100011001011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010100000111";
    r_D_in <= "0111000101011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010101010001001";
    r_D_in <= "0111111110010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100000111001000";
    r_D_in <= "0100110000111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111001001101";
    r_D_in <= "0110101110100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001010101010";
    r_D_in <= "0101101101010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100010001010";
    r_D_in <= "0111110000001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000001111000";
    r_D_in <= "0100101110101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111000110100";
    r_D_in <= "0100101001110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110101010101";
    r_D_in <= "0111000100010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010111000000";
    r_D_in <= "1001110001010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010001000010001";
    r_D_in <= "0101111101011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010111111100";
    r_D_in <= "0111101100010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100011110101101";
    r_D_in <= "0110010111110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101111010001";
    r_D_in <= "0110001101011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111110011001";
    r_D_in <= "0000110111011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011011011010";
    r_D_in <= "0111110010010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101000100110";
    r_D_in <= "0100101100010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100000100100000";
    r_D_in <= "0100001100110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100001100100";
    r_D_in <= "1001111100100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101110001001";
    r_D_in <= "0111010110111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111001011010";
    r_D_in <= "0110101000001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010011000010001";
    r_D_in <= "0011001010011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110000101011111";
    r_D_in <= "0110010101000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100110000001";
    r_D_in <= "0100100110010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111011111000";
    r_D_in <= "0101101001011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011010100010";
    r_D_in <= "0001101110100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000100011010";
    r_D_in <= "0010000101000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101110101111";
    r_D_in <= "0100110000100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111010010111";
    r_D_in <= "0100111011010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100001000110000";
    r_D_in <= "0111100101110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110011110001";
    r_D_in <= "0110101111001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011100010111";
    r_D_in <= "0101110000100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011000010010";
    r_D_in <= "1001110001011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111001101111";
    r_D_in <= "0111001010010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010101011011011";
    r_D_in <= "0101001011010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111110100110";
    r_D_in <= "0110110011001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110101111011010";
    r_D_in <= "0001101000110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000010011101";
    r_D_in <= "0101000011100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010111100111";
    r_D_in <= "0110011010001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011110000101";
    r_D_in <= "0110010000001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110001000111";
    r_D_in <= "0100001100111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111010110011";
    r_D_in <= "0011000101100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110010110110";
    r_D_in <= "0010100100110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000010011010";
    r_D_in <= "0101000011010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010100100010";
    r_D_in <= "0111000110010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100000110001";
    r_D_in <= "0110101000011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101010001101";
    r_D_in <= "1000111100011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111101010001";
    r_D_in <= "0010000011000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100010001010";
    r_D_in <= "0111101001100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100100010101";
    r_D_in <= "0001100000001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011101000111";
    r_D_in <= "1001111010010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101010001100000";
    r_D_in <= "0100001001101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100000010111";
    r_D_in <= "0111100111111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011100000111";
    r_D_in <= "0101110111100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010001001100";
    r_D_in <= "1001101110010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000101111001";
    r_D_in <= "0110111100110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100110100110";
    r_D_in <= "0111001001110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000111101001";
    r_D_in <= "0111010110010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011101000011";
    r_D_in <= "0101011110110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001111010110";
    r_D_in <= "0110100101110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010000001000";
    r_D_in <= "0111100110110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100000001100";
    r_D_in <= "0100111000011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001000101000001";
    r_D_in <= "1000011000110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110111011100";
    r_D_in <= "0101000001101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110111001111";
    r_D_in <= "0110101001000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010001110110";
    r_D_in <= "0101000010110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000000100010";
    r_D_in <= "0111111010000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011101101011";
    r_D_in <= "1010111101001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100011110000010";
    r_D_in <= "0111011011011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101100010101";
    r_D_in <= "0110110111011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110110000000";
    r_D_in <= "1010010101101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111001111000";
    r_D_in <= "0110001111011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010010101001";
    r_D_in <= "1001100011000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100110111111101";
    r_D_in <= "0111010000000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001100111101100";
    r_D_in <= "0100101100010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100100100100110";
    r_D_in <= "0101010111101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100111111101";
    r_D_in <= "0110001001000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100000110010";
    r_D_in <= "0110110111001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101000101001";
    r_D_in <= "0110100001001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110101111110101";
    r_D_in <= "0101101001111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011110010101";
    r_D_in <= "1000000011111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110010000010";
    r_D_in <= "1000111111001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101010011111";
    r_D_in <= "0111101010010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101101101011";
    r_D_in <= "0111110101100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011101101111";
    r_D_in <= "1000010000000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010001100000";
    r_D_in <= "1000000110100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011010000010";
    r_D_in <= "0101011110001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011001011000";
    r_D_in <= "0001011001000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110111111010";
    r_D_in <= "0110011011000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100111011111";
    r_D_in <= "0111000000011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110001100100";
    r_D_in <= "1001100101000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001001101100";
    r_D_in <= "1001010011000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110101111100010";
    r_D_in <= "0110110000011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000110011110";
    r_D_in <= "0110101101100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011011011011";
    r_D_in <= "1010101110011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101010010111001";
    r_D_in <= "0110101111010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100001001111111";
    r_D_in <= "0111001010111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111101001000";
    r_D_in <= "1000011100010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101010011000";
    r_D_in <= "0110111101010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110111100000";
    r_D_in <= "0111010011101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111100001001";
    r_D_in <= "1010011101100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011100000111";
    r_D_in <= "0111111000000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101110111100";
    r_D_in <= "0100000000000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110111101111";
    r_D_in <= "0100111101101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101100000000";
    r_D_in <= "0110110011111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010100000100";
    r_D_in <= "1000010000110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101101110100";
    r_D_in <= "0001101110111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101010011100100";
    r_D_in <= "0011110010001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010110100100";
    r_D_in <= "0101110111001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100000001000";
    r_D_in <= "0011101100100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011010001000";
    r_D_in <= "0101101100010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011100110010";
    r_D_in <= "0100110011010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011101100111";
    r_D_in <= "0101110010110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101100110110";
    r_D_in <= "0101000111010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100100011001011";
    r_D_in <= "0011111111100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101110011010111";
    r_D_in <= "0110111110010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010000000000";
    r_D_in <= "0101110101110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011011010001010";
    r_D_in <= "0011011010001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000100111101";
    r_D_in <= "0100001110111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011111010011";
    r_D_in <= "0111000000011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111110101000000";
    r_D_in <= "0000001100110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100101000010";
    r_D_in <= "0110101101110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001011100011010";
    r_D_in <= "0111001000010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100001110001";
    r_D_in <= "0101111010100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001100011100100";
    r_D_in <= "0110011110110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011001101110";
    r_D_in <= "0110011011011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011011100110";
    r_D_in <= "0111001010100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010101010000011";
    r_D_in <= "0110111100101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110101100011";
    r_D_in <= "0111101101010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111001010000";
    r_D_in <= "0100111010111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111011001000";
    r_D_in <= "0011101011010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011010110110";
    r_D_in <= "0111100101101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110010011110";
    r_D_in <= "0101001000000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111010001001";
    r_D_in <= "1000001111100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111100011101";
    r_D_in <= "0101011111101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110110101010";
    r_D_in <= "0100010110010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101100000100";
    r_D_in <= "0110110001100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001100000001";
    r_D_in <= "1010100010110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010100101010";
    r_D_in <= "0101001110010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101110110010100";
    r_D_in <= "0110011100001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110110111011";
    r_D_in <= "0101111011110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001100001011";
    r_D_in <= "0111100110100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010100110011";
    r_D_in <= "0010010110100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011100111000";
    r_D_in <= "1001010011000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101110000101";
    r_D_in <= "1000111110100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011000111100001";
    r_D_in <= "0110001110000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101010001110";
    r_D_in <= "0110000010101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010111111001";
    r_D_in <= "1000101000100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010011000010101";
    r_D_in <= "0100111000101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010010101000";
    r_D_in <= "0010111100101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010011110101000";
    r_D_in <= "0010011110101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010000011001";
    r_D_in <= "1000000101110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110100010001011";
    r_D_in <= "0111011010110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101101111010";
    r_D_in <= "0111110001001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100101101000";
    r_D_in <= "0111100000001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110000001010";
    r_D_in <= "0100110111100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101000100111";
    r_D_in <= "0111011001000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011001001010";
    r_D_in <= "1000010111000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101110000110001";
    r_D_in <= "0010111110001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111101101010";
    r_D_in <= "1000100101000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001001111100000";
    r_D_in <= "0011111100101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001100000110";
    r_D_in <= "0110100111010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001011101101101";
    r_D_in <= "0010011000001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111001011000111";
    r_D_in <= "0001011011100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010100011110";
    r_D_in <= "0011111111100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111010011000";
    r_D_in <= "1000000000001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010101000001100";
    r_D_in <= "0111010100110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010100010001";
    r_D_in <= "0011001000101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110010110011";
    r_D_in <= "0101011110000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101110101001";
    r_D_in <= "0111001110111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101010011101011";
    r_D_in <= "0011010010101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100100010000";
    r_D_in <= "1010010101000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010001110011";
    r_D_in <= "0101111011000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000000111100101";
    r_D_in <= "0111111010101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010100001111";
    r_D_in <= "1001111100011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000110000100100";
    r_D_in <= "0100110110010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111111000100";
    r_D_in <= "0011111110001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001010011100";
    r_D_in <= "0111111001010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110001000011";
    r_D_in <= "1000010011111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110111010000";
    r_D_in <= "0101111100000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111001100001";
    r_D_in <= "0111000010010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010110100110";
    r_D_in <= "0001110111111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000101100010";
    r_D_in <= "0010010000110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101001001110";
    r_D_in <= "0111101010001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100110100001";
    r_D_in <= "0110100111010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000000111101";
    r_D_in <= "0010001011101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101000001000011";
    r_D_in <= "0111100111101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000101110110";
    r_D_in <= "1000001010110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101101110101";
    r_D_in <= "0101100101110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110101001101";
    r_D_in <= "1000111000101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010111011111";
    r_D_in <= "0110011010110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011100011000";
    r_D_in <= "0101111100100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111101110000";
    r_D_in <= "0011010000110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111011011000";
    r_D_in <= "0110011000001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001000100101";
    r_D_in <= "1010000101110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000111110100";
    r_D_in <= "0011000011111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110101111101101";
    r_D_in <= "0110000100000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100110100000000";
    r_D_in <= "0100000101101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111111100110";
    r_D_in <= "0011010101101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010111110000";
    r_D_in <= "1010001001011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111110001001";
    r_D_in <= "0100100100110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110001110011";
    r_D_in <= "1000110110111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100001001100";
    r_D_in <= "0111100001001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100100011000";
    r_D_in <= "0001101110011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011000000001";
    r_D_in <= "0100101100110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110001100111011";
    r_D_in <= "0010100100110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101110011110";
    r_D_in <= "0000011111011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100000010000010";
    r_D_in <= "0110101001110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101010001110";
    r_D_in <= "0011111111011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001011110100110";
    r_D_in <= "1000000010001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001111000100";
    r_D_in <= "0111011100000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010001011101";
    r_D_in <= "1000010111101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110110110001";
    r_D_in <= "0100101001010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101110101100001";
    r_D_in <= "0101111111000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000011101011";
    r_D_in <= "0111111110110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111000001010010";
    r_D_in <= "0111011110100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101100110000011";
    r_D_in <= "1001101011010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110100100111";
    r_D_in <= "1001001000111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110001010111100";
    r_D_in <= "0111011110010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001001011011";
    r_D_in <= "1000000000010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100011001100";
    r_D_in <= "0110000010001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101111010111";
    r_D_in <= "0001111000010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000011010011";
    r_D_in <= "0101010001110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010011010010110";
    r_D_in <= "0110100011000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000101111101";
    r_D_in <= "0011101001010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101010011110";
    r_D_in <= "0100010011001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001010101000";
    r_D_in <= "1000011010111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111010101100";
    r_D_in <= "0001111011100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000010001000";
    r_D_in <= "0110000101110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101110100101";
    r_D_in <= "0010100011011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111000001100";
    r_D_in <= "1001100100101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001010101111111";
    r_D_in <= "0110110000010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111100001101";
    r_D_in <= "1000001100111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111010100111";
    r_D_in <= "0111111110001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010001101100101";
    r_D_in <= "0100111100100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111011110110";
    r_D_in <= "0011001110110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111100100000";
    r_D_in <= "0110101001101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100000110011";
    r_D_in <= "0111101101111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101010011001";
    r_D_in <= "0101110100101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100001101010";
    r_D_in <= "0110001110010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010110010000";
    r_D_in <= "0001110100110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111001000000";
    r_D_in <= "1000100100010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001100111111";
    r_D_in <= "1000011010111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000011110110";
    r_D_in <= "0110000011001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100000011001";
    r_D_in <= "0011001110011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110011000001";
    r_D_in <= "0101001110110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110101000100";
    r_D_in <= "1001101111001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101111000011";
    r_D_in <= "0111011111000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001011010101";
    r_D_in <= "0101010000110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010100011011";
    r_D_in <= "0111111111101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110000111000";
    r_D_in <= "0110011110001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010011001110101";
    r_D_in <= "0011111000010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010001000111111";
    r_D_in <= "0110000010101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010001011001";
    r_D_in <= "0111010111000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011110000000";
    r_D_in <= "1000010010000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010010000100";
    r_D_in <= "0110101000001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110101001010";
    r_D_in <= "0110111000010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011000100010";
    r_D_in <= "1001011011111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101010011001";
    r_D_in <= "0110000000001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110101101010001";
    r_D_in <= "0110111000110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111110100110";
    r_D_in <= "1000000010110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011000011011101";
    r_D_in <= "0110111000110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001101111111";
    r_D_in <= "0010110100001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111100111011";
    r_D_in <= "0111001110111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010100010010";
    r_D_in <= "0001010110001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001010111101";
    r_D_in <= "0100001100111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101110000111";
    r_D_in <= "0110000001111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001101111101";
    r_D_in <= "1000110010101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011100010010110";
    r_D_in <= "0110100000001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010111101010";
    r_D_in <= "1000001110000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011100000011";
    r_D_in <= "0110001110010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000110000111";
    r_D_in <= "0111101001001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110010011110";
    r_D_in <= "0111111100010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101101000100";
    r_D_in <= "0100110000011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000000101110011";
    r_D_in <= "0100001110011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001000110110111";
    r_D_in <= "0111110100101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111000000111";
    r_D_in <= "1000110011100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101101101010";
    r_D_in <= "0011101011001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000100100101";
    r_D_in <= "1000100010101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110010001111";
    r_D_in <= "0011000111110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001001100101110";
    r_D_in <= "0110100110101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110101111100001";
    r_D_in <= "0100000001110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100101000011";
    r_D_in <= "0011111100111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000110010100001";
    r_D_in <= "1000000111001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100000100100";
    r_D_in <= "1000001110100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111010001100";
    r_D_in <= "0011000101110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001100110110";
    r_D_in <= "0110111000101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010110010001";
    r_D_in <= "0110011000000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111111101000";
    r_D_in <= "0101100100001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110000111111110";
    r_D_in <= "1000001000001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111100111001";
    r_D_in <= "1011001010101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010100001011";
    r_D_in <= "0001100111011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111100100101";
    r_D_in <= "0100111100111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100110100100011";
    r_D_in <= "0100010101100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000000111110";
    r_D_in <= "0110011100000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010110011100";
    r_D_in <= "0111010111110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010101100100";
    r_D_in <= "0011111111001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011011101001";
    r_D_in <= "1010010101010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001010001101";
    r_D_in <= "0100110111111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110110110000100";
    r_D_in <= "0110110010110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010110111010";
    r_D_in <= "0001001011100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101000110010";
    r_D_in <= "0101001001001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010001111010";
    r_D_in <= "0111110101100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100101111101";
    r_D_in <= "0010000000011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101011010110";
    r_D_in <= "0100111010011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101110011111011";
    r_D_in <= "0101111001111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001101100010011";
    r_D_in <= "0110111110100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100010111100";
    r_D_in <= "0100111110011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010111111110";
    r_D_in <= "1000010111010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110011000011";
    r_D_in <= "0111010101100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001001010100";
    r_D_in <= "0100110110110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111000001011111";
    r_D_in <= "0111101010010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001111011100";
    r_D_in <= "0011001111110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111110101110110";
    r_D_in <= "0011110010011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010000011111";
    r_D_in <= "0100010101110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110101100001";
    r_D_in <= "0110110101100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101110100111110";
    r_D_in <= "1000101001100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111110011000";
    r_D_in <= "0111000110000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010001010001";
    r_D_in <= "0111011101101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011110000111";
    r_D_in <= "1001101100100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000011101000";
    r_D_in <= "0101001000011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001001100100010";
    r_D_in <= "0011010111101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010001110000";
    r_D_in <= "0111010100101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111111001011";
    r_D_in <= "0101111011000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010000101110";
    r_D_in <= "1001001010111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110100110101";
    r_D_in <= "1001001011111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110101010001";
    r_D_in <= "0011001111110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011101111110";
    r_D_in <= "0111011111111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001011000110010";
    r_D_in <= "0111010011010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110011101110";
    r_D_in <= "1011001000000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001001100010";
    r_D_in <= "1000001110000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110111101010";
    r_D_in <= "1000111111001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101110110110";
    r_D_in <= "0001011010001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110111111011";
    r_D_in <= "0110011110100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101111001001";
    r_D_in <= "0110101000100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000100101000110";
    r_D_in <= "0001000001100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001101110011";
    r_D_in <= "1010100001110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101010001111100";
    r_D_in <= "0111100111010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110100111100001";
    r_D_in <= "0110101111001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000010001011";
    r_D_in <= "0100000111000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001000101001";
    r_D_in <= "1000001101100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000101100101";
    r_D_in <= "0010100010010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101110001110101";
    r_D_in <= "0101110110101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111110000101";
    r_D_in <= "0011010000001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110001001111";
    r_D_in <= "0111110111010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111011011101";
    r_D_in <= "0010111101100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111110011011";
    r_D_in <= "1000010001010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101110110001";
    r_D_in <= "1000100001110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000011101111";
    r_D_in <= "0101100011010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000110000000011";
    r_D_in <= "1010110000111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101000111011";
    r_D_in <= "0111111011111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011110100101";
    r_D_in <= "0010100100011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100011011010";
    r_D_in <= "1001000001110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100110011000110";
    r_D_in <= "0100011001101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101001010001";
    r_D_in <= "0111000000000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100010000111";
    r_D_in <= "1001100010111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100010011110";
    r_D_in <= "0101111110011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101101001110";
    r_D_in <= "0101110100101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001101111000000";
    r_D_in <= "1010000001001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010010010101";
    r_D_in <= "0101110000010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110101111011";
    r_D_in <= "1001010111000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010110110101";
    r_D_in <= "0110011110001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110000011101";
    r_D_in <= "0011111001110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011110101011";
    r_D_in <= "1000011100000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100010001101";
    r_D_in <= "0001111101100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010101011110";
    r_D_in <= "0101010101101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010000111010";
    r_D_in <= "0101000111111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110101010100";
    r_D_in <= "0110010001000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110111010011";
    r_D_in <= "1010010011100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011111011010";
    r_D_in <= "0101100011111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000000011100111";
    r_D_in <= "0110111011101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011111101010";
    r_D_in <= "1000010001101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100000111000";
    r_D_in <= "0100011111110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101100110001";
    r_D_in <= "0110110001101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011000010001";
    r_D_in <= "0000101010010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000000001010";
    r_D_in <= "0111101101111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011100001110";
    r_D_in <= "1000110110110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101110001000";
    r_D_in <= "1000010011110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111100000001";
    r_D_in <= "1001111101110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110000101010";
    r_D_in <= "1000010011101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110010010000";
    r_D_in <= "1000010111100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001000010101";
    r_D_in <= "0111010000001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110111111000";
    r_D_in <= "0100110110110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110010000101";
    r_D_in <= "1000010110101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000011111100";
    r_D_in <= "0010111000000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000000111110100";
    r_D_in <= "0101110111110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010011010100101";
    r_D_in <= "0011001110000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111001110010";
    r_D_in <= "0100110100001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110011001010";
    r_D_in <= "1000011010111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010100110011";
    r_D_in <= "0100011101110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011010010011";
    r_D_in <= "1000110111000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011000111001001";
    r_D_in <= "0101011111010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001111001111110";
    r_D_in <= "0111010100001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100100000011";
    r_D_in <= "0101001010011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111010001110";
    r_D_in <= "0100111110000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010101001101111";
    r_D_in <= "0010111011001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001110011001";
    r_D_in <= "0111011101110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110110001001110";
    r_D_in <= "0111100001011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001011101000011";
    r_D_in <= "0011010101110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110001110110";
    r_D_in <= "0011110100110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100011000001001";
    r_D_in <= "1000110001010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111110011101";
    r_D_in <= "0110011000110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010101011101";
    r_D_in <= "0111100101111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011000000100";
    r_D_in <= "0101101100011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100010110001";
    r_D_in <= "0111110001000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101101110000";
    r_D_in <= "0110010110000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011101000110";
    r_D_in <= "1010010111101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100000000011";
    r_D_in <= "0101011111111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110000101011";
    r_D_in <= "0111001010111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110111001100";
    r_D_in <= "0100110111101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000110001100";
    r_D_in <= "0100110000100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001101010110";
    r_D_in <= "1001111111111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010100000111";
    r_D_in <= "0100101011111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100001000000";
    r_D_in <= "1001000011001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100010110011";
    r_D_in <= "0100111101100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110101010001111";
    r_D_in <= "0111000100100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111001001110010";
    r_D_in <= "0110110001100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111010010111";
    r_D_in <= "0111111001111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101101001110";
    r_D_in <= "0111100110111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100001001011";
    r_D_in <= "0111101000111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010111111000";
    r_D_in <= "0011100001010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010001101110";
    r_D_in <= "1010000101011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010101001010";
    r_D_in <= "0011011001011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110000111001011";
    r_D_in <= "1001001010010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110110001100";
    r_D_in <= "0010100110010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001101100101";
    r_D_in <= "0101110101100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000100000110011";
    r_D_in <= "0100101101010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111001101001";
    r_D_in <= "0101110110011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010100100010";
    r_D_in <= "0111000110100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101110101000";
    r_D_in <= "0110000101000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111110011010101";
    r_D_in <= "0111100101110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000110101111101";
    r_D_in <= "0011111101101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000101010100";
    r_D_in <= "0101001000110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001100111001";
    r_D_in <= "0100100010001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011101010101";
    r_D_in <= "0110011100001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001010001101101";
    r_D_in <= "0111110100100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110110000111";
    r_D_in <= "0010110010000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110001100101111";
    r_D_in <= "0110011011110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110000001111000";
    r_D_in <= "0111101111010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101000010100011";
    r_D_in <= "0011100010001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111011111111";
    r_D_in <= "0011111111010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001101010011";
    r_D_in <= "0100011010100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011000101000";
    r_D_in <= "1001010100100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000110000101";
    r_D_in <= "0101010010110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110010110110";
    r_D_in <= "0111000001111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000110010100101";
    r_D_in <= "0111010011101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111001010110";
    r_D_in <= "0011110011111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001000010101";
    r_D_in <= "0111001110011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010101010100";
    r_D_in <= "1000111011111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010100010001";
    r_D_in <= "0100000000100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011011110011";
    r_D_in <= "1000000011100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110110011110000";
    r_D_in <= "0101100001101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101110110000";
    r_D_in <= "0101100010000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101110011101";
    r_D_in <= "0111100010100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100100101100";
    r_D_in <= "0101101111101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011101101100";
    r_D_in <= "0011011111110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001001101010";
    r_D_in <= "0100110010110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010001100110";
    r_D_in <= "0100101100010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111101100001";
    r_D_in <= "1010001101010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111001111010101";
    r_D_in <= "0010000110100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011110001101";
    r_D_in <= "0001111000011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100101000111";
    r_D_in <= "0100010101101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110101011110";
    r_D_in <= "0110100101001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111010000101";
    r_D_in <= "0110100110100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001101100110";
    r_D_in <= "0101001110011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011000110011";
    r_D_in <= "1010110110111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100100110000";
    r_D_in <= "0110100100110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111000001010111";
    r_D_in <= "1001010111001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100010011001";
    r_D_in <= "1000011111111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101010101100000";
    r_D_in <= "0011101011000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010000010000";
    r_D_in <= "0101100011011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010111000010";
    r_D_in <= "0110010110110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100011011101";
    r_D_in <= "1001000010100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100010011011";
    r_D_in <= "0110111000010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010101110001";
    r_D_in <= "0011100100010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101110110110";
    r_D_in <= "1000011100010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101100011100001";
    r_D_in <= "0101111111000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100100100011";
    r_D_in <= "1010000010111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000100001000001";
    r_D_in <= "0101011111111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011011000010001";
    r_D_in <= "0100101101111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111011011110";
    r_D_in <= "0110001010000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111100010111";
    r_D_in <= "0100111100111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100010011101";
    r_D_in <= "0010111000101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110110111100";
    r_D_in <= "0011010010110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100011101001110";
    r_D_in <= "0101110100101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111010110101";
    r_D_in <= "1001100010001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011000111011";
    r_D_in <= "0110010110001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101111011010";
    r_D_in <= "0011011111100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000000110110100";
    r_D_in <= "0001010001100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000111011111110";
    r_D_in <= "1001000010101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001001110000";
    r_D_in <= "0101101101110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111001010000";
    r_D_in <= "0111001000110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110001110010011";
    r_D_in <= "0100000001111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110000100001";
    r_D_in <= "0111000000010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101110000000";
    r_D_in <= "1000100001001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100110010110001";
    r_D_in <= "0110000110100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001010110010";
    r_D_in <= "1000101100010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000000011100";
    r_D_in <= "0110001100101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110101101110001";
    r_D_in <= "1001100101001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001110101111";
    r_D_in <= "0101000111010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010000001001";
    r_D_in <= "0100100100111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110001111100010";
    r_D_in <= "0010010110100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110111000110";
    r_D_in <= "0011000110001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010001011111";
    r_D_in <= "0101010001111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010000010110";
    r_D_in <= "0101010010011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111000110100";
    r_D_in <= "0111111010010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111011101000";
    r_D_in <= "0010001010101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101111000110";
    r_D_in <= "0110001111000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101110111011010";
    r_D_in <= "0110000101000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010000101100";
    r_D_in <= "1000010100010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100100000011101";
    r_D_in <= "0011101011011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100001101011";
    r_D_in <= "0110011110010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111011100100";
    r_D_in <= "0101001110100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110000111110";
    r_D_in <= "0110001010110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111100010011";
    r_D_in <= "0101000011110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010001010100";
    r_D_in <= "0011110111100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100001011100100";
    r_D_in <= "0101010101100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010001110101001";
    r_D_in <= "1000000101010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110101110000011";
    r_D_in <= "1000100011001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010111001111";
    r_D_in <= "0110010111100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001001111100";
    r_D_in <= "0111101010000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001101110100";
    r_D_in <= "1000110011111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110001010011011";
    r_D_in <= "0111100110110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111100111100";
    r_D_in <= "1000111111101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101111100111";
    r_D_in <= "1000101010000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000000111100111";
    r_D_in <= "0001100100111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001101010000";
    r_D_in <= "0111000011010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011110010100";
    r_D_in <= "0101111110010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011000110000";
    r_D_in <= "0110111011101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001101011010";
    r_D_in <= "0111111100110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010110000100";
    r_D_in <= "1010001010011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100000111011";
    r_D_in <= "0010101001101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001110011000";
    r_D_in <= "0111111001001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010001011011";
    r_D_in <= "0110001110010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011110100111";
    r_D_in <= "0000111100000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101110110101";
    r_D_in <= "0010010111010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010000100011";
    r_D_in <= "0110010001000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100100011101";
    r_D_in <= "1000001011111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001010010010001";
    r_D_in <= "0111101111000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101110111110";
    r_D_in <= "0100101111110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110101101100111";
    r_D_in <= "0011101101100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101111101111";
    r_D_in <= "1000101000100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100001110010";
    r_D_in <= "1010010000110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001000010111";
    r_D_in <= "0111010000010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100001001000111";
    r_D_in <= "0100001010001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001110011110";
    r_D_in <= "1000001110011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100000001100";
    r_D_in <= "0111101111000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111000001101";
    r_D_in <= "0011100011101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101110111101";
    r_D_in <= "0101101010000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010101110100";
    r_D_in <= "1001110000001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010000010011";
    r_D_in <= "0100000101000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101110000000";
    r_D_in <= "0011100001010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101110000011010";
    r_D_in <= "1000010000110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000010010110";
    r_D_in <= "0100011010010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110110000111";
    r_D_in <= "1010010000001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010010010101";
    r_D_in <= "0110001111111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101001000101011";
    r_D_in <= "0101011111011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011100000001";
    r_D_in <= "0111000010001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110111111011";
    r_D_in <= "0110111001101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111001110000";
    r_D_in <= "0111101101110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101011111110";
    r_D_in <= "0011110100010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101101010111";
    r_D_in <= "0100101101101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000010010010";
    r_D_in <= "0110000011111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001111010101";
    r_D_in <= "0011010111011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010001101011";
    r_D_in <= "0111101101100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111100011110";
    r_D_in <= "0101001010010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111100100100";
    r_D_in <= "0100110000001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011110000101";
    r_D_in <= "0110010011001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011011111000";
    r_D_in <= "0001101110010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101111111101";
    r_D_in <= "0110111001100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011001000011";
    r_D_in <= "0110101000110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110000111111101";
    r_D_in <= "1000100000010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010111110010";
    r_D_in <= "0111111001101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010111110000";
    r_D_in <= "0110011011001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001000010111101";
    r_D_in <= "1001000110110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010011010111";
    r_D_in <= "0100000011101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001001000011";
    r_D_in <= "0101000110111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011101100001";
    r_D_in <= "0110010110011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011100001000011";
    r_D_in <= "0110111000110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101100101101111";
    r_D_in <= "0101110101111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010110101110";
    r_D_in <= "1000000010111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011111101011";
    r_D_in <= "0010011110000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101011100001";
    r_D_in <= "0111100010110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111110101101";
    r_D_in <= "0111100000110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101111110011";
    r_D_in <= "0100010100100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000011010000";
    r_D_in <= "1000000111011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101000110101011";
    r_D_in <= "0100100000111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011000110011";
    r_D_in <= "0100100101111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000010110011";
    r_D_in <= "0101101101000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111101100001";
    r_D_in <= "0101111101101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010011100011";
    r_D_in <= "0111011010101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001011101010";
    r_D_in <= "0000011011110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010011101001";
    r_D_in <= "0100111010100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011100100110011";
    r_D_in <= "0011101111000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010111000000";
    r_D_in <= "0011110101110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100011011101";
    r_D_in <= "0110000100101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101110000110";
    r_D_in <= "0010001110101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010011000100";
    r_D_in <= "1011000101000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110001111001";
    r_D_in <= "0011000001010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011000010011";
    r_D_in <= "1000100101001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111101110011";
    r_D_in <= "0010001101110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000110111001";
    r_D_in <= "0110001100011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111101111101";
    r_D_in <= "0101000011011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000100101000110";
    r_D_in <= "0110001100111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111010100000";
    r_D_in <= "0101110110111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001111010100011";
    r_D_in <= "0110010100110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001011100111";
    r_D_in <= "0100110000011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111010011011";
    r_D_in <= "0010001000100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100001110101101";
    r_D_in <= "1000110100011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010101011101";
    r_D_in <= "0111000100010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110100010111";
    r_D_in <= "0101101010101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011100011100";
    r_D_in <= "0111111010100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000111010000100";
    r_D_in <= "1000100111110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001011001010";
    r_D_in <= "0110110101101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010111100111";
    r_D_in <= "0100011110010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110100101110100";
    r_D_in <= "0111000101011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101000110101";
    r_D_in <= "0111011111010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101110001000001";
    r_D_in <= "0011111000100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010001111110";
    r_D_in <= "0001101110001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111100100000";
    r_D_in <= "0110111001100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101000010010";
    r_D_in <= "1000100110010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011001100000";
    r_D_in <= "0111111100110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101111010001";
    r_D_in <= "1010000110111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001101001011000";
    r_D_in <= "0110110011101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011001001001";
    r_D_in <= "1000011010100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100100111000";
    r_D_in <= "0101011000101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001101100010";
    r_D_in <= "1001110001001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110000001010101";
    r_D_in <= "0110110110010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000110011101000";
    r_D_in <= "0000110011101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001001001010001";
    r_D_in <= "0010000010010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101010101100";
    r_D_in <= "0011110010101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001101110110";
    r_D_in <= "0101100001101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001000110001";
    r_D_in <= "0101010110000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111100000010";
    r_D_in <= "0101110010101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100100111010";
    r_D_in <= "1000101011000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100000011010100";
    r_D_in <= "0100001000110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100001010010";
    r_D_in <= "0101101011101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000000101011101";
    r_D_in <= "0011110111011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011100001110";
    r_D_in <= "1000111101010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010110100100";
    r_D_in <= "0100101100000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011111000110";
    r_D_in <= "0000100111100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011100001011";
    r_D_in <= "0100101010011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101010101111100";
    r_D_in <= "0011100000101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011001110011";
    r_D_in <= "0110111100100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101100100010";
    r_D_in <= "0100001010111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011011000001";
    r_D_in <= "1001111111111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110100100001";
    r_D_in <= "0111111001010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110111010101";
    r_D_in <= "1000001010000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111001101110";
    r_D_in <= "0011111011010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001000001011010";
    r_D_in <= "1010100110001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011001110110";
    r_D_in <= "1001001101011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001111111111";
    r_D_in <= "1010011000011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001100001010100";
    r_D_in <= "0001100111000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000111110011100";
    r_D_in <= "1010001000011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111111010111";
    r_D_in <= "0111100001011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100001001110010";
    r_D_in <= "0100001100100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001110111010";
    r_D_in <= "0111100000101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101010000110";
    r_D_in <= "0100101101001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110000101011";
    r_D_in <= "0011111000011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101000111010";
    r_D_in <= "0110010101010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011101000001";
    r_D_in <= "0100110011100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000000010101000";
    r_D_in <= "1001010101101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001001111001000";
    r_D_in <= "0100001011011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000110110111011";
    r_D_in <= "0111001001100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101010100010";
    r_D_in <= "0111101011100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111000011111";
    r_D_in <= "0111111110110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010110101000";
    r_D_in <= "0101100001010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101000111011010";
    r_D_in <= "0100101001001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101110010001000";
    r_D_in <= "0110111010001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101011101001";
    r_D_in <= "1000111000100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010111101010";
    r_D_in <= "0101001001100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010100011011";
    r_D_in <= "0100000101111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110001001100010";
    r_D_in <= "1000000010000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011010010011";
    r_D_in <= "0111100110111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011001000000";
    r_D_in <= "1010001011101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011101001100";
    r_D_in <= "0110101010000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111000000101";
    r_D_in <= "0111110101010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000010000111";
    r_D_in <= "0110100000100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101110011010110";
    r_D_in <= "0111100100001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010001001101000";
    r_D_in <= "0011011101011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011010101001";
    r_D_in <= "0101100000101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010111010100";
    r_D_in <= "0011101001100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001011001001";
    r_D_in <= "0111010111110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010001011011";
    r_D_in <= "0100110101110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110000000000";
    r_D_in <= "0110111001100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111010100110";
    r_D_in <= "0101110010010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001011010111";
    r_D_in <= "0010101000010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101111001000";
    r_D_in <= "0100000101111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011110100100";
    r_D_in <= "0001011011011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110000110000";
    r_D_in <= "0110001010000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111111101100";
    r_D_in <= "0011100011011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110011110101";
    r_D_in <= "1000101000110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010101101110110";
    r_D_in <= "0011011101101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110111111011";
    r_D_in <= "0100011100001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000111100001110";
    r_D_in <= "1010011100111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111100000000";
    r_D_in <= "0111011000000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000110010011";
    r_D_in <= "0010000011110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101111101010";
    r_D_in <= "0001110011011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010010000101";
    r_D_in <= "0011110111110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100000000110000";
    r_D_in <= "0101001010000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001101000100100";
    r_D_in <= "0110111011101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010000111110";
    r_D_in <= "0011010010010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010001110011";
    r_D_in <= "0011010100010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101110110001";
    r_D_in <= "0110110111110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010100000011";
    r_D_in <= "0110010100111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101110000011";
    r_D_in <= "0111001000101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100110101110011";
    r_D_in <= "0011100100010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101001000001";
    r_D_in <= "0111110010001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100001010110";
    r_D_in <= "0101001011101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111110011110";
    r_D_in <= "0100111110100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101110000101110";
    r_D_in <= "0100111111100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010000010111";
    r_D_in <= "0010011110010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111111111111";
    r_D_in <= "0101000000000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101001001101";
    r_D_in <= "0001111100010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100011110011";
    r_D_in <= "1001000011111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010001001001110";
    r_D_in <= "0111111101001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010000111011";
    r_D_in <= "0101100111100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110111001101";
    r_D_in <= "0110010010001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010111101010";
    r_D_in <= "1000001101100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100111101100";
    r_D_in <= "0111100101100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101000000000";
    r_D_in <= "0111110111101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101001001111";
    r_D_in <= "0001000111111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111000101000";
    r_D_in <= "0110011000010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101001000001";
    r_D_in <= "0110001011001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100000011111";
    r_D_in <= "0101101010011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111110010110100";
    r_D_in <= "0100100001111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010011100110010";
    r_D_in <= "0110111100000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011100101101";
    r_D_in <= "0010100100001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111011100101";
    r_D_in <= "0110111000101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100111011100";
    r_D_in <= "0101100010101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000111111110";
    r_D_in <= "0011011001001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001000100000";
    r_D_in <= "0100011110101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000000011101";
    r_D_in <= "0111010100010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011001110100";
    r_D_in <= "1000111111101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011101001001";
    r_D_in <= "0100111000011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010011011000";
    r_D_in <= "1000110011111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100110010000";
    r_D_in <= "0010010101000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111011010100";
    r_D_in <= "0111100010000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111000001001";
    r_D_in <= "0100001110111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010110100110";
    r_D_in <= "1001001110101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001010011110111";
    r_D_in <= "0110101100110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110101111000";
    r_D_in <= "0100111111001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011000000010";
    r_D_in <= "0111101101101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111001101011";
    r_D_in <= "0111100111111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010011110011";
    r_D_in <= "0100001110011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111011000100";
    r_D_in <= "0001000011011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010110000101";
    r_D_in <= "0111001111001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010001111010";
    r_D_in <= "1010011001001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111111100111011";
    r_D_in <= "0000111010011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001100010010111";
    r_D_in <= "0101101110111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010101110111";
    r_D_in <= "0100011001000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111110010100";
    r_D_in <= "0100000100011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000011001011011";
    r_D_in <= "0111011100111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011011011011";
    r_D_in <= "0110011111001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011010111001";
    r_D_in <= "0110111011101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010110111000";
    r_D_in <= "0101011001000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001111100100110";
    r_D_in <= "0110000100010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111011000101";
    r_D_in <= "0011000010111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011010011101";
    r_D_in <= "1000010111101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111001110111";
    r_D_in <= "0111111101111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101110101000111";
    r_D_in <= "0101111100000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010010101111100";
    r_D_in <= "0100110001000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110110101011111";
    r_D_in <= "0100111010111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001110010001";
    r_D_in <= "0100000110110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001010010010100";
    r_D_in <= "1010011011010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111111101110";
    r_D_in <= "0110000000001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010001000111001";
    r_D_in <= "0111001100100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111001011100";
    r_D_in <= "1000010010001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001010010001";
    r_D_in <= "1000000000001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011011100110101";
    r_D_in <= "0110111101000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110010101100101";
    r_D_in <= "0111000011000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010001101011001";
    r_D_in <= "0110000010000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001111000011";
    r_D_in <= "0101000100011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100100110101";
    r_D_in <= "0111000111001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001111010100011";
    r_D_in <= "0100110001110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001010111110011";
    r_D_in <= "0111110000000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111101101100";
    r_D_in <= "1000011101101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111011011001110";
    r_D_in <= "0111011101010000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100101101011";
    r_D_in <= "0110010010111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100010111110";
    r_D_in <= "0101001001000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000010010100000";
    r_D_in <= "1000001110011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110100001110";
    r_D_in <= "0101111010111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011011001100110";
    r_D_in <= "0101101010010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010101001110";
    r_D_in <= "1000111011110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101100000011";
    r_D_in <= "0101100000100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110100111010";
    r_D_in <= "0100100110011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010110011110";
    r_D_in <= "0101001010100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100010000100";
    r_D_in <= "0001111011001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110111010010";
    r_D_in <= "0101101101111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111010111101";
    r_D_in <= "0001110011000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000101011110";
    r_D_in <= "0110101100101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100111001011";
    r_D_in <= "0001101011001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011011100101";
    r_D_in <= "1001101000000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100000010111011";
    r_D_in <= "0100000011101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111110000110";
    r_D_in <= "1000000101000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010111101111";
    r_D_in <= "0100000111100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000000111101011";
    r_D_in <= "0101011011101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110111010010100";
    r_D_in <= "0110111011100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011010011101";
    r_D_in <= "0111111110010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110101001111111";
    r_D_in <= "0010111010100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110101101111";
    r_D_in <= "0011100100011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100101101011";
    r_D_in <= "0101011011000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101100100111";
    r_D_in <= "0101110111100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101110101100";
    r_D_in <= "0011100100101100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010010000111011";
    r_D_in <= "0101110110010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100111011101";
    r_D_in <= "1000111100001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111101111100";
    r_D_in <= "0101000011000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010100101011";
    r_D_in <= "0010011111110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001001110100";
    r_D_in <= "1001010000111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110000111001000";
    r_D_in <= "0110101010010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110111100100";
    r_D_in <= "0111111000001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111101000111";
    r_D_in <= "1001011011000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011000110100000";
    r_D_in <= "0100111010110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001101001110011";
    r_D_in <= "0010000000010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010001010101111";
    r_D_in <= "0111111100100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001101111111";
    r_D_in <= "0000010010110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100100011111010";
    r_D_in <= "0100101000111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111000111111";
    r_D_in <= "0110010101111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110110001001";
    r_D_in <= "0101100001100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111110100101";
    r_D_in <= "0101100000100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000001100100101";
    r_D_in <= "1001101111110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110101001100";
    r_D_in <= "0111111100000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111111010001";
    r_D_in <= "0001001001000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111111011101";
    r_D_in <= "0110011100101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100100001110100";
    r_D_in <= "0101101100110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001011010011";
    r_D_in <= "1000011000100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001111100101";
    r_D_in <= "0110100001101110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000000110001010";
    r_D_in <= "0111000101111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100000010000";
    r_D_in <= "1000111010110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001100011101";
    r_D_in <= "0110011110011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010110100000";
    r_D_in <= "0110101001001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100100100110000";
    r_D_in <= "0011110000110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000010110111";
    r_D_in <= "0101011000110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110000110110010";
    r_D_in <= "0110010100100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101110011000111";
    r_D_in <= "0101110011001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111100001110";
    r_D_in <= "1000001000100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111110100100";
    r_D_in <= "0111101000100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010100100011100";
    r_D_in <= "0111010101001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010101101001";
    r_D_in <= "0111011011000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011100011000011";
    r_D_in <= "0101001110111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001111101001011";
    r_D_in <= "0110101100011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111001100000001";
    r_D_in <= "0001100101011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000000100101100";
    r_D_in <= "0000001001011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100110101100010";
    r_D_in <= "0101100011110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000001101011111";
    r_D_in <= "0000100001111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110001111111010";
    r_D_in <= "0110010000110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011011100010";
    r_D_in <= "0100111111001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101000101000";
    r_D_in <= "0111011001000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011111010100";
    r_D_in <= "0010001110011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100010010000";
    r_D_in <= "0101111101110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010100001010";
    r_D_in <= "0110100111010010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100011110110001";
    r_D_in <= "0110110010111111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000110100100111";
    r_D_in <= "0111001110000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010010010010";
    r_D_in <= "1001011111010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110101101000";
    r_D_in <= "0101010011111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111101001001110";
    r_D_in <= "1010001011101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110101111101001";
    r_D_in <= "0010111001010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001111001010";
    r_D_in <= "0111001010101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001000010011100";
    r_D_in <= "1000100111010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111110111000011";
    r_D_in <= "0001011011000010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001010101101001";
    r_D_in <= "0100000110011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111001110011";
    r_D_in <= "0111110101011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100110101000001";
    r_D_in <= "0101000111000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100110011100";
    r_D_in <= "0011111010111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111011011010";
    r_D_in <= "1001011011001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000010101010";
    r_D_in <= "0101101100001100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101000100110";
    r_D_in <= "0100000001001110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101011101000000";
    r_D_in <= "0010101110011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111100101110";
    r_D_in <= "0110100011010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111100110110110";
    r_D_in <= "1000011011000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101100011101101";
    r_D_in <= "0101100011110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001001110010110";
    r_D_in <= "0100010011011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111101011100";
    r_D_in <= "0101011101101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010111011111";
    r_D_in <= "0101011000000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111010110110101";
    r_D_in <= "1001110100101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100010111001";
    r_D_in <= "1001111110101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110011000101010";
    r_D_in <= "0110101000111110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011010011110";
    r_D_in <= "0110110011110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100000001111";
    r_D_in <= "0101100000011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001101000000011";
    r_D_in <= "0111010101111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101110001010";
    r_D_in <= "0011010010011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101011110001";
    r_D_in <= "0011111000101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001111000100000";
    r_D_in <= "0111001110110001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000110001010110";
    r_D_in <= "0111101100101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110000100000";
    r_D_in <= "0110100000011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000011110101";
    r_D_in <= "0111001110100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000111100100111";
    r_D_in <= "1000100000001010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111100011100";
    r_D_in <= "0110111110100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010000010100011";
    r_D_in <= "0101111110101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100110100010111";
    r_D_in <= "0101101001011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010111001011000";
    r_D_in <= "0101101101100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101110110111000";
    r_D_in <= "0010001011001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011001010001011";
    r_D_in <= "0110011000010110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010110010101101";
    r_D_in <= "0101100111011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010011010101100";
    r_D_in <= "0011001010001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111011010100";
    r_D_in <= "0001111011110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010111010100111";
    r_D_in <= "0011111001011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101111001110110";
    r_D_in <= "0010100000100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011000011010001";
    r_D_in <= "0011100001000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011100101111";
    r_D_in <= "1000100110111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100111101111";
    r_D_in <= "0100100111101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101110000011000";
    r_D_in <= "0110111110100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101010001101";
    r_D_in <= "1001000011010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101011000100";
    r_D_in <= "0111011100011100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000100110100";
    r_D_in <= "0111010111100011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111111010011";
    r_D_in <= "0110001110001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010011010000101";
    r_D_in <= "0010110000101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011101000000101";
    r_D_in <= "1000100101101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110110000000100";
    r_D_in <= "0100110000011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000110111010101";
    r_D_in <= "0010110101100001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010100001100";
    r_D_in <= "0101100010001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101010101001";
    r_D_in <= "0101110001101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010001100110";
    r_D_in <= "0100111101110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011110110010100";
    r_D_in <= "1000100111011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111110100010111";
    r_D_in <= "1000000000001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010010000101";
    r_D_in <= "0100101010101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001101011100011";
    r_D_in <= "0110100010011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011100001010001";
    r_D_in <= "0101101100100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101101011001100";
    r_D_in <= "0110001000100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111001000100101";
    r_D_in <= "1001010111011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110011000101101";
    r_D_in <= "1001111110010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011111101000110";
    r_D_in <= "0110001010101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111101110110";
    r_D_in <= "0001011000110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101000111000110";
    r_D_in <= "0101110110111000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011010000000";
    r_D_in <= "0111011011001000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010100001110101";
    r_D_in <= "0100111101011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100001111110";
    r_D_in <= "0100101101011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001110011101001";
    r_D_in <= "0111111010011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001000110110010";
    r_D_in <= "0101001111110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101011100101";
    r_D_in <= "0100001111011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101100001101100";
    r_D_in <= "0111100111011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100011101000101";
    r_D_in <= "0101101100010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111100111000";
    r_D_in <= "0110010011011011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100011101110101";
    r_D_in <= "0011100010001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001011000110011";
    r_D_in <= "1010010001010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110111100010000";
    r_D_in <= "0101000110010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100001100011";
    r_D_in <= "0111011010011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011010110111110";
    r_D_in <= "0110100000101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010001111001010";
    r_D_in <= "0110010101111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010101110110011";
    r_D_in <= "0010110101011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111000101100";
    r_D_in <= "0010000100011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101111010000111";
    r_D_in <= "0110000010100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100010101000001";
    r_D_in <= "0111011011000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101000000111111";
    r_D_in <= "0100011101011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110110010111111";
    r_D_in <= "1000010101111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110111001100";
    r_D_in <= "0101010110101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001010100110110";
    r_D_in <= "0111101101111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100111101000010";
    r_D_in <= "0110100011101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000111101110100";
    r_D_in <= "1000010110001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100011110100";
    r_D_in <= "1001001011001011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001101101000100";
    r_D_in <= "0110111100011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010101110101111";
    r_D_in <= "0111100000000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100101101000001";
    r_D_in <= "0011110111110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101001111010";
    r_D_in <= "0111010100100111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100001000010";
    r_D_in <= "0111111000010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001011100011001";
    r_D_in <= "0111001110110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010001011111100";
    r_D_in <= "0111000100000100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010011100111100";
    r_D_in <= "0111101000000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101001100001001";
    r_D_in <= "1000011011001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110000100101100";
    r_D_in <= "0010111010110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000111100000";
    r_D_in <= "0111111001100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010010110001";
    r_D_in <= "0111011100100110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000101000100";
    r_D_in <= "0010100100010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100110100100100";
    r_D_in <= "0111000010011001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000011000011000";
    r_D_in <= "0111100111101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111000001111000";
    r_D_in <= "0111000001111010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0001110101000001";
    r_D_in <= "0101110000100000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101011110000101";
    r_D_in <= "0110011100101101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111011011011101";
    r_D_in <= "0100000000000000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001011111001";
    r_D_in <= "0100110110101111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101111011011";
    r_D_in <= "0111000110010100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111001011101010";
    r_D_in <= "0111100010110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001111011100";
    r_D_in <= "1000110110011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110001001101110";
    r_D_in <= "0100111011111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110000011110100";
    r_D_in <= "0110100010110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110100000010111";
    r_D_in <= "0100110110000011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111100010010010";
    r_D_in <= "0100111001011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011010000000010";
    r_D_in <= "0101110100110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100011011101";
    r_D_in <= "0111000100110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111010011110";
    r_D_in <= "0101100110110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000111111111";
    r_D_in <= "0110001001111011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100101011001101";
    r_D_in <= "0110101001110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011001001011101";
    r_D_in <= "1000110010101011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011100000011011";
    r_D_in <= "1000100000100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000010111010000";
    r_D_in <= "0101001000110011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011110010000101";
    r_D_in <= "0100111101100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0110100110100110";
    r_D_in <= "0111111001100100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1011111100111000";
    r_D_in <= "0100000011111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001100010101000";
    r_D_in <= "0110111111100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000111011001100";
    r_D_in <= "0010010010110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001001000101110";
    r_D_in <= "1000100010010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000101101101";
    r_D_in <= "0111100011110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010101010001011";
    r_D_in <= "1000001101111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110011101011";
    r_D_in <= "0101110001110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000110001000100";
    r_D_in <= "0111010000110000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111000000110001";
    r_D_in <= "0000111111010111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101111000111";
    r_D_in <= "1000000011010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011011111011010";
    r_D_in <= "0110100100111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1001011010001101";
    r_D_in <= "0110111100000110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111111010101011";
    r_D_in <= "1000100000000001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111000010001101";
    r_D_in <= "1000100111010101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101000000000101";
    r_D_in <= "0011000011001101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0011101111011010";
    r_D_in <= "1000001011010011";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010011100110";
    r_D_in <= "0010111001001001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010110001000010";
    r_D_in <= "0010110110110111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101000010110101";
    r_D_in <= "0100101110100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111110000001000";
    r_D_in <= "0010110101000101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111101110011";
    r_D_in <= "0110010011111101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100010011110010";
    r_D_in <= "0100010011111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101010000010000";
    r_D_in <= "1000001011110110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1100000111010111";
    r_D_in <= "0011111110110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000110100100010";
    r_D_in <= "1010001110001111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100111000010101";
    r_D_in <= "1001010111011110";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1101010100000100";
    r_D_in <= "0011000011011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000100011100000";
    r_D_in <= "1001001111111001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110010111100011";
    r_D_in <= "0001111110101001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1000101110110101";
    r_D_in <= "0111010101000111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101011010001";
    r_D_in <= "0110011001011101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1010101111010100";
    r_D_in <= "0111000000110100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0111000100110000";
    r_D_in <= "0111110010011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000000001100101";
    r_D_in <= "0010110001111100";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111110000000110";
    r_D_in <= "0100100110101010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010000010110110";
    r_D_in <= "0100100001110101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111101110000000";
    r_D_in <= "0111001111011111";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1111010011101010";
    r_D_in <= "0100101101100101";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101011111101";
    r_D_in <= "0010101000110010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0010001110001100";
    r_D_in <= "0010010110010001";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0101101001100100";
    r_D_in <= "0111000101011010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "1110110010001110";
    r_D_in <= "0101000001101000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0000101111000101";
    r_D_in <= "0111000010011000";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;
    r_N_in <= "0100001011001100";
    r_D_in <= "0100011011100010";
    output_tmp := to_integer(signed(w_Q_out));
    WRITE (line_out, output_tmp);
    WRITELINE(file_out, line_out);
    wait for 10 ns;


  end process;
  
End Behavioral;