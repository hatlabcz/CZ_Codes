library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity test_integrator_tb is	
end test_integrator_tb;

architecture Behavioral of test_integrator_tb is
  
  constant r_input_width : integer:=16;
  constant c_clk_period  : time:=10 ns;
 
  
  signal r_ch1_data0       : std_logic_vector(r_input_width-1 downto 0); -- Signal
  signal r_ch1_data1       : std_logic_vector(r_input_width-1 downto 0); -- Signal
  signal r_ch1_data2       : std_logic_vector(r_input_width-1 downto 0); -- Signal
  signal r_ch1_data3       : std_logic_vector(r_input_width-1 downto 0); -- Signal
  signal r_ch1_data4       : std_logic_vector(r_input_width-1 downto 0); -- Signal
  signal r_ch1_valid       : std_logic := '1'; -- Signal
  
  signal SI : std_logic_vector(31 downto 0);
  signal SQ : std_logic_vector(31 downto 0);
  signal RI : std_logic_vector(31 downto 0);
  signal RQ : std_logic_vector(31 downto 0);

  
  signal r_rst     : std_logic:='0';
  signal r_clk     : std_logic:='0';
 
 
  component Integrator_v1 is	
	Generic (
		input_width : integer := 16;
		output_width : integer := 32;
		input_signed : boolean := TRUE;
		input_latch	: boolean := TRUE;
		points : integer := 10
	);
	Port (
		Din_sdi_dataStreamFCx5_S_data_0 : in std_logic_vector(input_width-1 downto 0);
		Din_sdi_dataStreamFCx5_S_data_1 : in std_logic_vector(input_width-1 downto 0);
		Din_sdi_dataStreamFCx5_S_data_2 : in std_logic_vector(input_width-1 downto 0);
		Din_sdi_dataStreamFCx5_S_data_3 : in std_logic_vector(input_width-1 downto 0);
		Din_sdi_dataStreamFCx5_S_data_4 : in std_logic_vector(input_width-1 downto 0);
		Din_sdi_dataStreamFCx5_S_valid : in std_logic;
		
		
		Dout : out std_logic_vector(output_width-1 downto 0);
		
		clk : in std_logic;
		rst : in std_logic;
		clr : in std_logic
	);
  end component Integrator_v1;
  

begin

  p_clk_gen : process is
    begin 
	  wait for c_clk_period/2;
	  r_clk <= not(r_clk);
  end process p_clk_gen;
  
  Integrator_1 : Integrator_v1
    port map (
      rst     => r_rst,
	  clr     => r_rst,
	  clk     => r_clk,
	  
      Din_sdi_dataStreamFCx5_S_data_0  => r_ch1_data0,
	  Din_sdi_dataStreamFCx5_S_data_1  => r_ch1_data1,
	  Din_sdi_dataStreamFCx5_S_data_2  => r_ch1_data2,
	  Din_sdi_dataStreamFCx5_S_data_3  => r_ch1_data3,
	  Din_sdi_dataStreamFCx5_S_data_4  => r_ch1_data4,
	  Din_sdi_dataStreamFCx5_S_valid   => r_ch1_valid,
	 
	  Dout => SI
      );
	  

  process
  begin
    
        r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "1111111111111111";
    r_ch1_data2 <= "1111111111111111";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000001";
    r_ch1_data1 <= "0000000000000001";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111111111111111";
    wait for 10 ns;
    r_ch1_data0 <= "1111111111111111";
    r_ch1_data1 <= "1111111111111111";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000001";
    r_ch1_data4 <= "0000000000000010";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000001";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111111111111111";
    r_ch1_data3 <= "1111111111111110";
    r_ch1_data4 <= "1111111111111110";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000001";
    r_ch1_data2 <= "0000000000000011";
    r_ch1_data3 <= "0000000000000011";
    r_ch1_data4 <= "0000000000000010";
    wait for 10 ns;
    r_ch1_data0 <= "1111111111111110";
    r_ch1_data1 <= "1111111111111100";
    r_ch1_data2 <= "1111111111111100";
    r_ch1_data3 <= "1111111111111110";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000101";
    r_ch1_data1 <= "0000000000000101";
    r_ch1_data2 <= "0000000000000011";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111111111111101";
    wait for 10 ns;
    r_ch1_data0 <= "1111111111111010";
    r_ch1_data1 <= "1111111111111100";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000100";
    r_ch1_data4 <= "0000000000000111";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000101";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111111111111011";
    r_ch1_data3 <= "1111111111110111";
    r_ch1_data4 <= "1111111111110111";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000110";
    r_ch1_data2 <= "0000000000001011";
    r_ch1_data3 <= "0000000000001011";
    r_ch1_data4 <= "0000000000000111";
    wait for 10 ns;
    r_ch1_data0 <= "1111111111111000";
    r_ch1_data1 <= "1111111111110011";
    r_ch1_data2 <= "1111111111110010";
    r_ch1_data3 <= "1111111111110111";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000010000";
    r_ch1_data1 <= "0000000000010001";
    r_ch1_data2 <= "0000000000001011";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111111111110100";
    wait for 10 ns;
    r_ch1_data0 <= "1111111111101011";
    r_ch1_data1 <= "1111111111110011";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000001110";
    r_ch1_data4 <= "0000000000011000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000010000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111111111101111";
    r_ch1_data3 <= "1111111111100011";
    r_ch1_data4 <= "1111111111100010";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000010101";
    r_ch1_data2 <= "0000000000100011";
    r_ch1_data3 <= "0000000000100101";
    r_ch1_data4 <= "0000000000010111";
    wait for 10 ns;
    r_ch1_data0 <= "1111111111100111";
    r_ch1_data1 <= "1111111111010110";
    r_ch1_data2 <= "1111111111010100";
    r_ch1_data3 <= "1111111111100100";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000110011";
    r_ch1_data1 <= "0000000000110101";
    r_ch1_data2 <= "0000000000100010";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111111111011100";
    wait for 10 ns;
    r_ch1_data0 <= "1111111111000001";
    r_ch1_data1 <= "1111111111011000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000101011";
    r_ch1_data4 <= "0000000001001001";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000110000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111111111001101";
    r_ch1_data3 <= "1111111110101010";
    r_ch1_data4 <= "1111111110100111";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000111101";
    r_ch1_data2 <= "0000000001100111";
    r_ch1_data3 <= "0000000001101010";
    r_ch1_data4 <= "0000000001000100";
    wait for 10 ns;
    r_ch1_data0 <= "1111111110111000";
    r_ch1_data1 <= "1111111110000111";
    r_ch1_data2 <= "1111111110000011";
    r_ch1_data3 <= "1111111110110000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000010001111";
    r_ch1_data1 <= "0000000010010100";
    r_ch1_data2 <= "0000000001011110";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111111110011011";
    wait for 10 ns;
    r_ch1_data0 <= "1111111101010010";
    r_ch1_data1 <= "1111111110010001";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000001110110";
    r_ch1_data4 <= "0000000011000110";
    wait for 10 ns;
    r_ch1_data0 <= "0000000010000010";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111111101110101";
    r_ch1_data3 <= "1111111100011000";
    r_ch1_data4 <= "1111111100010001";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000010100010";
    r_ch1_data2 <= "0000000100001111";
    r_ch1_data3 <= "0000000100010111";
    r_ch1_data4 <= "0000000010110010";
    wait for 10 ns;
    r_ch1_data0 <= "1111111101000011";
    r_ch1_data1 <= "1111111011000100";
    r_ch1_data2 <= "1111111010111011";
    r_ch1_data3 <= "1111111100110001";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000101101111";
    r_ch1_data1 <= "0000000101111010";
    r_ch1_data2 <= "0000000011110001";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111111100000001";
    wait for 10 ns;
    r_ch1_data0 <= "1111111001001010";
    r_ch1_data1 <= "1111111011101001";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000100100111";
    r_ch1_data4 <= "0000000111101100";
    wait for 10 ns;
    r_ch1_data0 <= "0000000101000010";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111111010101011";
    r_ch1_data3 <= "1111110111001000";
    r_ch1_data4 <= "1111110110111000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000110001000";
    r_ch1_data2 <= "0000001010001101";
    r_ch1_data3 <= "0000001010100000";
    r_ch1_data4 <= "0000000110101011";
    wait for 10 ns;
    r_ch1_data0 <= "1111111000111101";
    r_ch1_data1 <= "1111110100010010";
    r_ch1_data2 <= "1111110011111101";
    r_ch1_data3 <= "1111111000010111";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000001101011011";
    r_ch1_data1 <= "0000001101110010";
    r_ch1_data2 <= "0000001000110000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111110110110010";
    wait for 10 ns;
    r_ch1_data0 <= "1111110000010001";
    r_ch1_data1 <= "1111110110000010";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000001010100000";
    r_ch1_data4 <= "0000010001011101";
    wait for 10 ns;
    r_ch1_data0 <= "0000001011010111";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111110100000011";
    r_ch1_data3 <= "1111101100001011";
    r_ch1_data4 <= "1111101011101010";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000001101100011";
    r_ch1_data2 <= "0000010110011111";
    r_ch1_data3 <= "0000010111000011";
    r_ch1_data4 <= "0000001110100110";
    wait for 10 ns;
    r_ch1_data0 <= "1111110000101011";
    r_ch1_data1 <= "1111100110100101";
    r_ch1_data2 <= "1111100101111101";
    r_ch1_data3 <= "1111101111100001";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000011100101010";
    r_ch1_data1 <= "0000011101010111";
    r_ch1_data2 <= "0000010010100101";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111101100100010";
    wait for 10 ns;
    r_ch1_data0 <= "1111011111000000";
    r_ch1_data1 <= "1111101011001000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000010101110111";
    r_ch1_data4 <= "0000100100001100";
    wait for 10 ns;
    r_ch1_data0 <= "0000010111011010";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111100111100001";
    r_ch1_data3 <= "1111010111100000";
    r_ch1_data4 <= "1111010110100101";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000011011010110";
    r_ch1_data2 <= "0000101101001111";
    r_ch1_data3 <= "0000101110001110";
    r_ch1_data4 <= "0000011101001100";
    wait for 10 ns;
    r_ch1_data0 <= "1111100001100010";
    r_ch1_data1 <= "1111001101101000";
    r_ch1_data2 <= "1111001100100011";
    r_ch1_data3 <= "1111011111100001";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000110111111110";
    r_ch1_data1 <= "0000111001001001";
    r_ch1_data2 <= "0000100100000011";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111011010011100";
    wait for 10 ns;
    r_ch1_data0 <= "1111000000101101";
    r_ch1_data1 <= "1111011000000110";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000101001100011";
    r_ch1_data4 <= "0001000100100100";
    wait for 10 ns;
    r_ch1_data0 <= "0000101100000101";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111010010001011";
    r_ch1_data3 <= "1110110100011001";
    r_ch1_data4 <= "1110110010111011";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000110010011100";
    r_ch1_data2 <= "0001010011001011";
    r_ch1_data3 <= "0001010100101111";
    r_ch1_data4 <= "0000110101010111";
    wait for 10 ns;
    r_ch1_data0 <= "1111001000101001";
    r_ch1_data1 <= "1110100100110000";
    r_ch1_data2 <= "1110100011000101";
    r_ch1_data3 <= "1111000101100001";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0001100011110111";
    r_ch1_data1 <= "0001100101101010";
    r_ch1_data2 <= "0000111111111100";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1110111101110010";
    wait for 10 ns;
    r_ch1_data0 <= "1110010001000101";
    r_ch1_data1 <= "1110111010010001";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0001001000001010";
    r_ch1_data4 <= "0001110110101111";
    wait for 10 ns;
    r_ch1_data0 <= "0001001011111000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1110110001100110";
    r_ch1_data3 <= "1101111111000010";
    r_ch1_data4 <= "1101111100111011";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0001010101000001";
    r_ch1_data2 <= "0010001011110000";
    r_ch1_data3 <= "0010001101111110";
    r_ch1_data4 <= "0001011001001000";
    wait for 10 ns;
    r_ch1_data0 <= "1110100100000101";
    r_ch1_data1 <= "1101101000111101";
    r_ch1_data2 <= "1101100110101000";
    r_ch1_data3 <= "1110011111110001";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0010100010110111";
    r_ch1_data1 <= "0010100101010010";
    r_ch1_data2 <= "0001100111101010";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1110010101010011";
    wait for 10 ns;
    r_ch1_data0 <= "1101001110010110";
    r_ch1_data1 <= "1110010000101001";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0001110010100010";
    r_ch1_data4 <= "0010111011111001";
    wait for 10 ns;
    r_ch1_data0 <= "0001110111010110";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1110000101011001";
    r_ch1_data3 <= "1100110110111100";
    r_ch1_data4 <= "1100110100010000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0010000010111101";
    r_ch1_data2 <= "0011010110101000";
    r_ch1_data3 <= "0011011001011000";
    r_ch1_data4 <= "0010001000000011";
    wait for 10 ns;
    r_ch1_data0 <= "1101110100100000";
    r_ch1_data1 <= "1100011011011111";
    r_ch1_data2 <= "1100011000101010";
    r_ch1_data3 <= "1101101111010010";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0011110010101110";
    r_ch1_data1 <= "0011110101100101";
    r_ch1_data2 <= "0010011001100011";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1101100010111000";
    wait for 10 ns;
    r_ch1_data0 <= "1011111011111101";
    r_ch1_data1 <= "1101011101011111";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0010100110001001";
    r_ch1_data4 <= "0100001111110000";
    wait for 10 ns;
    r_ch1_data0 <= "0010101011100101";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1101010000110010";
    r_ch1_data3 <= "1011100001100010";
    r_ch1_data4 <= "1011011110100101";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0010111000010110";
    r_ch1_data2 <= "0100101101001111";
    r_ch1_data3 <= "0100110000001100";
    r_ch1_data4 <= "0010111101110100";
    wait for 10 ns;
    r_ch1_data0 <= "1100111110100011";
    r_ch1_data1 <= "1011000100000010";
    r_ch1_data2 <= "1011000001000110";
    r_ch1_data3 <= "1100111001000110";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0101001010100110";
    r_ch1_data1 <= "0101001101100000";
    r_ch1_data2 <= "0011001111111010";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1100101100100010";
    wait for 10 ns;
    r_ch1_data0 <= "1010100100000111";
    r_ch1_data1 <= "1100100111001111";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0011011100010001";
    r_ch1_data4 <= "0101100111001101";
    wait for 10 ns;
    r_ch1_data0 <= "0011100001011100";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1100011011001010";
    r_ch1_data3 <= "1010001010111110";
    r_ch1_data4 <= "1010001000010001";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0011101101001011";
    r_ch1_data2 <= "0110000010011010";
    r_ch1_data3 <= "0110000101000010";
    r_ch1_data4 <= "0011110010000010";
    wait for 10 ns;
    r_ch1_data0 <= "1100001010110011";
    r_ch1_data1 <= "1001110000101111";
    r_ch1_data2 <= "1001101110001110";
    r_ch1_data3 <= "1100000110001010";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0110011011100010";
    r_ch1_data1 <= "0110011101111010";
    r_ch1_data2 <= "0100000001010000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1011111011111010";
    wait for 10 ns;
    r_ch1_data0 <= "1001010110101010";
    r_ch1_data1 <= "1011110111110001";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0100001010111001";
    r_ch1_data4 <= "0110110001111100";
    wait for 10 ns;
    r_ch1_data0 <= "0100001110101110";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1011101110110110";
    r_ch1_data3 <= "1001000100000101";
    r_ch1_data4 <= "1001000010001100";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0100010110111001";
    r_ch1_data2 <= "0111000101000000";
    r_ch1_data3 <= "0111000110101101";
    r_ch1_data4 <= "0100011010000011";
    wait for 10 ns;
    r_ch1_data0 <= "1011100011111110";
    r_ch1_data1 <= "1000110010111001";
    r_ch1_data2 <= "1000110001011001";
    r_ch1_data3 <= "1011100001001100";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0111010100001101";
    r_ch1_data1 <= "0111010101011111";
    r_ch1_data2 <= "0100100010111011";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1011011011100111";
    wait for 10 ns;
    r_ch1_data0 <= "1000100100101110";
    r_ch1_data1 <= "1011011001101001";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0100100111100011";
    r_ch1_data4 <= "0111011111000110";
    wait for 10 ns;
    r_ch1_data0 <= "0100101001000111";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1011010110000000";
    r_ch1_data3 <= "1000011101001011";
    r_ch1_data4 <= "1000011100100101";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0100101011101110";
    r_ch1_data2 <= "0111100101010111";
    r_ch1_data3 <= "0111100101101111";
    r_ch1_data4 <= "0100101100011001";
    wait for 10 ns;
    r_ch1_data0 <= "1011010011010100";
    r_ch1_data1 <= "1000011001010011";
    r_ch1_data2 <= "1000011001001011";
    r_ch1_data3 <= "1011010011000110";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0111100110110101";
    r_ch1_data1 <= "0111100110101101";
    r_ch1_data2 <= "0100101100101100";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1011010011100111";
    wait for 10 ns;
    r_ch1_data0 <= "1000011010101001";
    r_ch1_data1 <= "1011010100010010";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0100101011000111";
    r_ch1_data4 <= "0111100011011011";
    wait for 10 ns;
    r_ch1_data0 <= "0100101010000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1011010110111001";
    r_ch1_data3 <= "1000100000000100";
    r_ch1_data4 <= "1000100000111010";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0100100110010111";
    r_ch1_data2 <= "0111011011010010";
    r_ch1_data3 <= "0111011010001101";
    r_ch1_data4 <= "0100100100011001";
    wait for 10 ns;
    r_ch1_data0 <= "1011011101000101";
    r_ch1_data1 <= "1000101010100001";
    r_ch1_data2 <= "1000101011110011";
    r_ch1_data3 <= "1011011111011110";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0111001110100111";
    r_ch1_data1 <= "0111001101000111";
    r_ch1_data2 <= "0100011100000010";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1011100101111101";
    wait for 10 ns;
    r_ch1_data0 <= "1000111011000000";
    r_ch1_data1 <= "1011101001000111";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0100010100101011";
    r_ch1_data4 <= "0110111101110100";
    wait for 10 ns;
    r_ch1_data0 <= "0100010001001010";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1011110001010010";
    r_ch1_data3 <= "1001001100000000";
    r_ch1_data4 <= "1001001110000100";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0100001000001111";
    r_ch1_data2 <= "0110101001010110";
    r_ch1_data3 <= "0110100111000111";
    r_ch1_data4 <= "0100000100000110";
    wait for 10 ns;
    r_ch1_data0 <= "1011111110110000";
    r_ch1_data1 <= "1001100010000110";
    r_ch1_data2 <= "1001100100011110";
    r_ch1_data3 <= "1100000011001001";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0110010001110010";
    r_ch1_data1 <= "0110001111010001";
    r_ch1_data2 <= "0011110101001101";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1100001101111110";
    wait for 10 ns;
    r_ch1_data0 <= "1001111101100110";
    r_ch1_data1 <= "1100010010110101";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0011101001111000";
    r_ch1_data4 <= "0101110111101111";
    wait for 10 ns;
    r_ch1_data0 <= "0011100100110110";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1100011110100100";
    r_ch1_data3 <= "1010010110000000";
    r_ch1_data4 <= "1010011000110011";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0011011000110001";
    r_ch1_data2 <= "0101011011111001";
    r_ch1_data3 <= "0101011001000010";
    r_ch1_data4 <= "0011010011011110";
    wait for 10 ns;
    r_ch1_data0 <= "1100110000000110";
    r_ch1_data1 <= "1010110010100000";
    r_ch1_data2 <= "1010110101011010";
    r_ch1_data3 <= "1100110101011111";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0100111110111010";
    r_ch1_data1 <= "0100111011111110";
    r_ch1_data2 <= "0011000001011101";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1101000010001100";
    wait for 10 ns;
    r_ch1_data0 <= "1011010010110001";
    r_ch1_data1 <= "1101000111101010";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0010110100101100";
    r_ch1_data4 <= "0100100001011011";
    wait for 10 ns;
    r_ch1_data0 <= "0010101111001110";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1101010100011011";
    r_ch1_data3 <= "1011101101010100";
    r_ch1_data4 <= "1011110000010000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0010100010100001";
    r_ch1_data2 <= "0100000100000011";
    r_ch1_data3 <= "0100000001001001";
    r_ch1_data4 <= "0010011101001000";
    wait for 10 ns;
    r_ch1_data0 <= "1101100110011101";
    r_ch1_data1 <= "1100001010011011";
    r_ch1_data2 <= "1100001101010010";
    r_ch1_data3 <= "1101101011110001";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0011100111010110";
    r_ch1_data1 <= "0011100100100001";
    r_ch1_data2 <= "0010001011100000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1101110111111101";
    wait for 10 ns;
    r_ch1_data0 <= "1100101001011000";
    r_ch1_data1 <= "1101111101000011";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0001111111100101";
    r_ch1_data4 <= "0011001011110000";
    wait for 10 ns;
    r_ch1_data0 <= "0001111010100111";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1110001000101010";
    r_ch1_data3 <= "1101000001100000";
    r_ch1_data4 <= "1101000100000111";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0001101111010111";
    r_ch1_data2 <= "0010110001101010";
    r_ch1_data3 <= "0010101111001001";
    r_ch1_data4 <= "0001101010101101";
    wait for 10 ns;
    r_ch1_data0 <= "1110011000010110";
    r_ch1_data1 <= "1101011010101110";
    r_ch1_data2 <= "1101011101001001";
    r_ch1_data3 <= "1110011100110110";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0010011001011000";
    r_ch1_data1 <= "0010010111000011";
    r_ch1_data2 <= "0001011011111011";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1110100110111000";
    wait for 10 ns;
    r_ch1_data0 <= "1101110100010000";
    r_ch1_data1 <= "1110101010111111";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0001010010010101";
    r_ch1_data4 <= "0010000011000101";
    wait for 10 ns;
    r_ch1_data0 <= "0001001110011010";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1110110100001000";
    r_ch1_data3 <= "1110000111010001";
    r_ch1_data4 <= "1110001001010001";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0001000101101111";
    r_ch1_data2 <= "0001101110111011";
    r_ch1_data3 <= "0001101101000010";
    r_ch1_data4 <= "0001000010001110";
    wait for 10 ns;
    r_ch1_data0 <= "1111000000000100";
    r_ch1_data1 <= "1110011010010110";
    r_ch1_data2 <= "1110011100001001";
    r_ch1_data3 <= "1111000011011000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0001011100111011";
    r_ch1_data1 <= "0001011011010000";
    r_ch1_data2 <= "0000110111010111";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111001010101001";
    wait for 10 ns;
    r_ch1_data0 <= "1110101100110101";
    r_ch1_data1 <= "1111001101100100";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000110000100011";
    r_ch1_data4 <= "0001001101000101";
    wait for 10 ns;
    r_ch1_data0 <= "0000101101110101";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111010011111011";
    r_ch1_data3 <= "1110111010000100";
    r_ch1_data4 <= "1110111011011100";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000100111111010";
    r_ch1_data2 <= "0000111111010011";
    r_ch1_data3 <= "0000111110000010";
    r_ch1_data4 <= "0000100101100100";
    wait for 10 ns;
    r_ch1_data0 <= "1111011011111101";
    r_ch1_data1 <= "1111000110110111";
    r_ch1_data2 <= "1111001000000010";
    r_ch1_data3 <= "1111011110001000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000110011011101";
    r_ch1_data1 <= "0000110010011000";
    r_ch1_data2 <= "0000011110011110";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111100010110100";
    wait for 10 ns;
    r_ch1_data0 <= "1111010010110001";
    r_ch1_data1 <= "1111100100101010";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000011010001011";
    r_ch1_data4 <= "0000101001011011";
    wait for 10 ns;
    r_ch1_data0 <= "0000011000011111";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111101000100110";
    r_ch1_data3 <= "1111011010111111";
    r_ch1_data4 <= "1111011011110100";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000010100111000";
    r_ch1_data2 <= "0000100001000000";
    r_ch1_data3 <= "0000100000010000";
    r_ch1_data4 <= "0000010011011110";
    wait for 10 ns;
    r_ch1_data0 <= "1111101101011011";
    r_ch1_data1 <= "1111100010101001";
    r_ch1_data2 <= "1111100011010110";
    r_ch1_data3 <= "1111101110101101";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000011010000011";
    r_ch1_data1 <= "0000011001011011";
    r_ch1_data2 <= "0000001111010101";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111110001011010";
    wait for 10 ns;
    r_ch1_data0 <= "1111101001100001";
    r_ch1_data1 <= "1111110010011101";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000001100111001";
    r_ch1_data4 <= "0000010100010110";
    wait for 10 ns;
    r_ch1_data0 <= "0000001011111101";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111110100101001";
    r_ch1_data3 <= "1111101110000110";
    r_ch1_data4 <= "1111101110100011";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000001001111110";
    r_ch1_data2 <= "0000001111101111";
    r_ch1_data3 <= "0000001111010100";
    r_ch1_data4 <= "0000001001001110";
    wait for 10 ns;
    r_ch1_data0 <= "1111110111010000";
    r_ch1_data1 <= "1111110010001110";
    r_ch1_data2 <= "1111110010100101";
    r_ch1_data3 <= "1111110111111100";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000001100000011";
    r_ch1_data1 <= "0000001011101110";
    r_ch1_data2 <= "0000000111000011";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111111001010101";
    wait for 10 ns;
    r_ch1_data0 <= "1111110101110011";
    r_ch1_data1 <= "1111111001111000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000101110011";
    r_ch1_data4 <= "0000001001001000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000101010101";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111111010111110";
    r_ch1_data3 <= "1111111000000101";
    r_ch1_data4 <= "1111111000010100";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000100010111";
    r_ch1_data2 <= "0000000110110110";
    r_ch1_data3 <= "0000000110101010";
    r_ch1_data4 <= "0000000011111111";
    wait for 10 ns;
    r_ch1_data0 <= "1111111100001111";
    r_ch1_data1 <= "1111111010000110";
    r_ch1_data2 <= "1111111010010001";
    r_ch1_data3 <= "1111111100100100";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000101000101";
    r_ch1_data1 <= "0000000100111100";
    r_ch1_data2 <= "0000000010111101";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111111101001110";
    wait for 10 ns;
    r_ch1_data0 <= "1111111011110001";
    r_ch1_data1 <= "1111111101011110";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000010011000";
    r_ch1_data4 <= "0000000011101111";
    wait for 10 ns;
    r_ch1_data0 <= "0000000010001011";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111111101111110";
    r_ch1_data3 <= "1111111100110100";
    r_ch1_data4 <= "1111111100111010";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000001101111";
    r_ch1_data2 <= "0000000010101110";
    r_ch1_data3 <= "0000000010101001";
    r_ch1_data4 <= "0000000001100101";
    wait for 10 ns;
    r_ch1_data0 <= "1111111110100010";
    r_ch1_data1 <= "1111111101101100";
    r_ch1_data2 <= "1111111101110001";
    r_ch1_data3 <= "1111111110101011";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000001111101";
    r_ch1_data1 <= "0000000001111001";
    r_ch1_data2 <= "0000000001001000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111111110111100";
    wait for 10 ns;
    r_ch1_data0 <= "1111111110011001";
    r_ch1_data1 <= "1111111111000011";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000111001";
    r_ch1_data4 <= "0000000001011001";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000110011";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111111111010000";
    r_ch1_data3 <= "1111111110110101";
    r_ch1_data4 <= "1111111110110111";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000101000";
    r_ch1_data2 <= "0000000000111111";
    r_ch1_data3 <= "0000000000111101";
    r_ch1_data4 <= "0000000000100100";
    wait for 10 ns;
    r_ch1_data0 <= "1111111111011110";
    r_ch1_data1 <= "1111111111001011";
    r_ch1_data2 <= "1111111111001101";
    r_ch1_data3 <= "1111111111100010";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000101100";
    r_ch1_data1 <= "0000000000101010";
    r_ch1_data2 <= "0000000000011001";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111111111101001";
    wait for 10 ns;
    r_ch1_data0 <= "1111111111011101";
    r_ch1_data1 <= "1111111111101011";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000010011";
    r_ch1_data4 <= "0000000000011110";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000010001";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111111111110000";
    r_ch1_data3 <= "1111111111100111";
    r_ch1_data4 <= "1111111111101000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000001101";
    r_ch1_data2 <= "0000000000010101";
    r_ch1_data3 <= "0000000000010100";
    r_ch1_data4 <= "0000000000001100";
    wait for 10 ns;
    r_ch1_data0 <= "1111111111110101";
    r_ch1_data1 <= "1111111111101111";
    r_ch1_data2 <= "1111111111110000";
    r_ch1_data3 <= "1111111111110111";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000001110";
    r_ch1_data1 <= "0000000000001101";
    r_ch1_data2 <= "0000000000001000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111111111111001";
    wait for 10 ns;
    r_ch1_data0 <= "1111111111110101";
    r_ch1_data1 <= "1111111111111010";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000110";
    r_ch1_data4 <= "0000000000001001";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000101";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111111111111011";
    r_ch1_data3 <= "1111111111111001";
    r_ch1_data4 <= "1111111111111001";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000100";
    r_ch1_data2 <= "0000000000000110";
    r_ch1_data3 <= "0000000000000110";
    r_ch1_data4 <= "0000000000000011";
    wait for 10 ns;
    r_ch1_data0 <= "1111111111111101";
    r_ch1_data1 <= "1111111111111011";
    r_ch1_data2 <= "1111111111111011";
    r_ch1_data3 <= "1111111111111110";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000100";
    r_ch1_data1 <= "0000000000000100";
    r_ch1_data2 <= "0000000000000010";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "1111111111111110";
    wait for 10 ns;
    r_ch1_data0 <= "1111111111111101";
    r_ch1_data1 <= "1111111111111111";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000001";
    r_ch1_data4 <= "0000000000000010";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000001";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "1111111111111111";
    r_ch1_data3 <= "1111111111111110";
    r_ch1_data4 <= "1111111111111110";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000001";
    r_ch1_data2 <= "0000000000000001";
    r_ch1_data3 <= "0000000000000001";
    r_ch1_data4 <= "0000000000000001";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "1111111111111111";
    r_ch1_data2 <= "1111111111111111";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000001";
    r_ch1_data1 <= "0000000000000001";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";
    r_ch1_data3 <= "0000000000000000";
    r_ch1_data4 <= "0000000000000000";
    wait for 10 ns;
    r_ch1_data0 <= "0000000000000000";
    r_ch1_data1 <= "0000000000000000";
    r_ch1_data2 <= "0000000000000000";

  
  end process;
  
End Behavioral;